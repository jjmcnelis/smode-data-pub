9c9
< 		time:units = "days since 1950-01-01T00:00:00" ;
---
> 		time:units = "days since 1950-01-01 00:00:00" ;
12c12
< 		longitude:_FillValue = NaN ;
---
> 		longitude::_FillValue = -9999. ;
16d15
< 		longitude:axis = "X" ;
19c18
< 		longitude:coverage_content_type = "coordinate" ;
---
> 		longitude:coverage_content_type = "referenceInformation" ;
21c20
< 		latitude:_FillValue = NaN ;
---
> 		latitude::_FillValue = -9999. ;
25d23
< 		latitude:axis = "Y" ;
28c26
< 		latitude:coverage_content_type = "coordinate" ;
---
> 		latitude:coverage_content_type = "referenceInformation" ;
30c28
< 		sst:_FillValue = NaN ;
---
> 		sst::_FillValue = -9999. ;
41c39
< 		sss:_FillValue = NaN ;
---
> 		sss::_FillValue = -9999. ;
52c50
< 		solar_radiation:_FillValue = NaN ;
---
> 		solar_radiation::_FillValue = -9999. ;
63c61
< 		long_radiation:_FillValue = NaN ;
---
> 		long_radiation::_FillValue = -9999. ;
74c72
< 		pressure:_FillValue = NaN ;
---
> 		pressure::_FillValue = -9999. ;
85c83
< 		wind_direction:_FillValue = NaN ;
---
> 		wind_direction::_FillValue = -9999. ;
97c95
< 		wind_speed_5m:_FillValue = NaN ;
---
> 		wind_speed_5m::_FillValue = -9999. ;
108c106
< 		relative_humidity_2m:_FillValue = NaN ;
---
> 		relative_humidity_2m::_FillValue = -9999. ;
119c117
< 		specific_humidity_2m:_FillValue = NaN ;
---
> 		specific_humidity_2m::_FillValue = -9999. ;
130c128
< 		air_temperature_2m:_FillValue = NaN ;
---
> 		air_temperature_2m::_FillValue = -9999. ;
141c139
< 		wind_speed_10m:_FillValue = NaN ;
---
> 		wind_speed_10m::_FillValue = -9999. ;
152c150
< 		relative_humidity_10m:_FillValue = NaN ;
---
> 		relative_humidity_10m::_FillValue = -9999. ;
163c161
< 		specific_humidity_10m:_FillValue = NaN ;
---
> 		specific_humidity_10m::_FillValue = -9999. ;
174c172
< 		air_temperature_10m:_FillValue = NaN ;
---
> 		air_temperature_10m::_FillValue = -9999. ;
192c190
< 		:id = "PO.DAAC-SMODE-SDRON" ;
---
> 		:id = "PODAAC-SMODE-SDRON" ;
197c195
< 		:source = "TBD" ;
---
> 		:source = "S-MODE_PFC_saildrone_##.nc.cdl" ;
226,227c224,225
< 		:geospatial_lat_units = "degrees" ;
< 		:geospatial_lat_resolution = "0.1" ;
---
> 		:geospatial_lat_units = "degrees_north" ;
> 		:geospatial_lat_resolution = "0.1 degrees" ;
230,231c228,229
< 		:geospatial_lon_units = "degrees" ;
< 		:geospatial_lon_resolution = "0.1" ;
---
> 		:geospatial_lon_units = "degrees_east" ;
> 		:geospatial_lon_resolution = "0.1 degrees" ;
234,235c232,233
< 		:geospatial_vertical_resolution = "1" ;
< 		:geospatial_vertical_units = "m" ;
---
> 		:geospatial_vertical_resolution = "1 meters" ;
> 		:geospatial_vertical_units = "meters" ;
237,239c235,237
< 		:time_coverage_start = "16-Oct-2017" ;
< 		:time_coverage_end = "17-Nov-2017" ;
< 		:date_created = "01-Sep-2020 14:13:03" ;
---
> 		:time_coverage_start = "2017-11-16THH:MM:SS" ;
> 		:time_coverage_end = "2017-11-17HH:MM:SS" ;
> 		:date_created = "2020-09-01T14:13:03" ;
