netcdf S-MODE_PFC_OC2004B_meteorology_\#\# {
dimensions:
	time = 43200 ;
variables:
	double time(time) ;
		time:long_name = "Time" ;
		time:comment = "Time from Ships Data Files" ;
		time:axis = "T" ;
		time:standard_name = "time" ;
		time:units = "days since 1950-01-01 00:00:00" ;
		time:coverage_content_type = "coordinate" ;
	double latitude(time) ;
		latitude:_FillValue = -9999. ;
		latitude:long_name = "Latitude" ;
		latitude:comment = "Latitude from Ships Data Files" ;
		latitude:valid_max = 90. ;
		latitude:valid_min = -90. ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "referenceInformation" ;
	double longitude(time) ;
		longitude:_FillValue = -9999. ;
		longitude:long_name = "Longitude" ;
		longitude:comment = "Longitude from Ships Data Files" ;
		longitude:valid_max = 180. ;
		longitude:valid_min = -180. ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "referenceInformation" ;
	double speed_over_ground(time) ;
		speed_over_ground:_FillValue = -9999. ;
		speed_over_ground:long_name = "Speed Over Ground from Ships Data Files" ;
		speed_over_ground:valid_max = 7.01995752416612 ;
		speed_over_ground:valid_min = 0.00121450605039624 ;
		speed_over_ground:add_offset = 0. ;
		speed_over_ground:scale_factor = 1. ;
		speed_over_ground:standard_name = "platform_speed_wrt_ground" ;
		speed_over_ground:units = "m s-1" ;
		speed_over_ground:coverage_content_type = "physicalMeasurement" ;
		speed_over_ground:coordinates = "time longitude latitude" ;
	double course_over_ground(time) ;
		course_over_ground:_FillValue = -9999. ;
		course_over_ground:long_name = "Course Over Ground from Ships Data Files" ;
		course_over_ground:valid_max = 360. ;
		course_over_ground:valid_min = 0. ;
		course_over_ground:add_offset = 0. ;
		course_over_ground:scale_factor = 1. ;
		course_over_ground:standard_name = "platform_course" ;
		course_over_ground:units = "degrees" ;
		course_over_ground:coverage_content_type = "physicalMeasurement" ;
		course_over_ground:coordinates = "time longitude latitude" ;
	double heading(time) ;
		heading:_FillValue = -9999. ;
		heading:long_name = "Heading from Ships Data Files" ;
		heading:valid_max = 360. ;
		heading:valid_min = 0. ;
		heading:add_offset = 0. ;
		heading:scale_factor = 1. ;
		heading:standard_name = "heading" ;
		heading:units = "degrees" ;
		heading:coverage_content_type = "physicalMeasurement" ;
		heading:coordinates = "time longitude latitude" ;
	double eastward_current(time) ;
		eastward_current:_FillValue = -9999. ;
		eastward_current:long_name = "Eastward Current from ADCP Measurement" ;
		eastward_current:valid_max = 2. ;
		eastward_current:valid_min = -2. ;
		eastward_current:add_offset = 0. ;
		eastward_current:scale_factor = 1. ;
		eastward_current:standard_name = "eastward_sea_water_velocity" ;
		eastward_current:units = "m s-1" ;
		eastward_current:coverage_content_type = "physicalMeasurement" ;
		eastward_current:coordinates = "time longitude latitude" ;
	double northward_current(time) ;
		northward_current:_FillValue = -9999. ;
		northward_current:long_name = "Northward Current from ADCP Measurement" ;
		northward_current:valid_max = 2. ;
		northward_current:valid_min = -2. ;
		northward_current:add_offset = 0. ;
		northward_current:scale_factor = 1. ;
		northward_current:standard_name = "northward_sea_water_velocity" ;
		northward_current:units = "m s-1" ;
		northward_current:coverage_content_type = "physicalMeasurement" ;
		northward_current:coordinates = "time longitude latitude" ;
	double wind_speed_relative_to_earth_18m(time) ;
		wind_speed_relative_to_earth_18m:_FillValue = -9999. ;
		wind_speed_relative_to_earth_18m:long_name = "Wind Speed relative to Earth at ~18m from Sonic Anemometers on the bow mast" ;
		wind_speed_relative_to_earth_18m:valid_max = 13.6921813602126 ;
		wind_speed_relative_to_earth_18m:valid_min = 0. ;
		wind_speed_relative_to_earth_18m:add_offset = 0. ;
		wind_speed_relative_to_earth_18m:scale_factor = 1. ;
		wind_speed_relative_to_earth_18m:standard_name = "wind_speed" ;
		wind_speed_relative_to_earth_18m:units = "m s-1" ;
		wind_speed_relative_to_earth_18m:coverage_content_type = "physicalMeasurement" ;
		wind_speed_relative_to_earth_18m:coordinates = "time longitude latitude" ;
	double wind_direction_relative_to_earth(time) ;
		wind_direction_relative_to_earth:_FillValue = -9999. ;
		wind_direction_relative_to_earth:long_name = "Wind Direction relative to Earth from Sonic Anemometers on the bow mast" ;
		wind_direction_relative_to_earth:valid_max = 360. ;
		wind_direction_relative_to_earth:valid_min = 0. ;
		wind_direction_relative_to_earth:add_offset = 0. ;
		wind_direction_relative_to_earth:scale_factor = 1. ;
		wind_direction_relative_to_earth:standard_name = "wind_from_direction" ;
		wind_direction_relative_to_earth:units = "degrees" ;
		wind_direction_relative_to_earth:coverage_content_type = "physicalMeasurement" ;
		wind_direction_relative_to_earth:coordinates = "time longitude latitude" ;
	double wind_speed_relative_to_earth(time) ;
		wind_speed_relative_to_earth:_FillValue = -9999. ;
		wind_speed_relative_to_earth:long_name = "Wind Speed relative to Earth adjusted to 10m computed from ADCP measurements" ;
		wind_speed_relative_to_earth:valid_max = 13.0163613641973 ;
		wind_speed_relative_to_earth:valid_min = 0. ;
		wind_speed_relative_to_earth:add_offset = 0. ;
		wind_speed_relative_to_earth:scale_factor = 1. ;
		wind_speed_relative_to_earth:standard_name = "wind_speed" ;
		wind_speed_relative_to_earth:units = "m s-1" ;
		wind_speed_relative_to_earth:coverage_content_type = "physicalMeasurement" ;
		wind_speed_relative_to_earth:coordinates = "time longitude latitude" ;
	double neutral_wind_speed_relative_to_earth(time) ;
		neutral_wind_speed_relative_to_earth:_FillValue = -9999. ;
		neutral_wind_speed_relative_to_earth:long_name = "Neutral Wind Speed relative to Earth adjusted to 10m and neutral stratification computed from ADCP measurements" ;
		neutral_wind_speed_relative_to_earth:valid_max = 13.1644591886842 ;
		neutral_wind_speed_relative_to_earth:valid_min = 0. ;
		neutral_wind_speed_relative_to_earth:add_offset = 0. ;
		neutral_wind_speed_relative_to_earth:scale_factor = 1. ;
		neutral_wind_speed_relative_to_earth:standard_name = "wind_speed" ;
		neutral_wind_speed_relative_to_earth:units = "m s-1" ;
		neutral_wind_speed_relative_to_earth:coverage_content_type = "physicalMeasurement" ;
		neutral_wind_speed_relative_to_earth:coordinates = "time longitude latitude" ;
	double wind_speed_relative_to_water_18m(time) ;
		wind_speed_relative_to_water_18m:_FillValue = -9999. ;
		wind_speed_relative_to_water_18m:long_name = "Wind Speed relative to water at ~18m from Sonic Anemometers on the bow mast" ;
		wind_speed_relative_to_water_18m:valid_max = 13.7852907180786 ;
		wind_speed_relative_to_water_18m:valid_min = 0. ;
		wind_speed_relative_to_water_18m:add_offset = 0. ;
		wind_speed_relative_to_water_18m:scale_factor = 1. ;
		wind_speed_relative_to_water_18m:standard_name = "wind_speed" ;
		wind_speed_relative_to_water_18m:units = "m s-1" ;
		wind_speed_relative_to_water_18m:coverage_content_type = "physicalMeasurement" ;
		wind_speed_relative_to_water_18m:coordinates = "time longitude latitude" ;
	double wind_direction_relative_to_water(time) ;
		wind_direction_relative_to_water:_FillValue = -9999. ;
		wind_direction_relative_to_water:long_name = "Wind Direction relative to water from Sonic Anemometers on the bow mast" ;
		wind_direction_relative_to_water:valid_max = 360. ;
		wind_direction_relative_to_water:valid_min = 0. ;
		wind_direction_relative_to_water:add_offset = 0. ;
		wind_direction_relative_to_water:scale_factor = 1. ;
		wind_direction_relative_to_water:standard_name = "wind_from_direction" ;
		wind_direction_relative_to_water:units = "degrees" ;
		wind_direction_relative_to_water:coverage_content_type = "physicalMeasurement" ;
		wind_direction_relative_to_water:coordinates = "time longitude latitude" ;
	double wind_speed_relative_to_water_2m(time) ;
		wind_speed_relative_to_water_2m:_FillValue = -9999. ;
		wind_speed_relative_to_water_2m:long_name = "Wind Speed relative to water adjusted to 2m computed from ADCP measurements" ;
		wind_speed_relative_to_water_2m:valid_max = 11.1033296585083 ;
		wind_speed_relative_to_water_2m:valid_min = 0. ;
		wind_speed_relative_to_water_2m:add_offset = 0. ;
		wind_speed_relative_to_water_2m:scale_factor = 1. ;
		wind_speed_relative_to_water_2m:standard_name = "wind_speed" ;
		wind_speed_relative_to_water_2m:units = "m s-1" ;
		wind_speed_relative_to_water_2m:coverage_content_type = "physicalMeasurement" ;
		wind_speed_relative_to_water_2m:coordinates = "time longitude latitude" ;
	double wind_speed_relative_to_water_10m(time) ;
		wind_speed_relative_to_water_10m:_FillValue = -9999. ;
		wind_speed_relative_to_water_10m:long_name = "Wind Speed relative to water adjusted to 10m computed from ADCP measurements" ;
		wind_speed_relative_to_water_10m:valid_max = 13.1284875869751 ;
		wind_speed_relative_to_water_10m:valid_min = 0. ;
		wind_speed_relative_to_water_10m:add_offset = 0. ;
		wind_speed_relative_to_water_10m:scale_factor = 1. ;
		wind_speed_relative_to_water_10m:standard_name = "wind_speed" ;
		wind_speed_relative_to_water_10m:units = "m s-1" ;
		wind_speed_relative_to_water_10m:coverage_content_type = "physicalMeasurement" ;
		wind_speed_relative_to_water_10m:coordinates = "time longitude latitude" ;
	double neutral_wind_speed_relative_to_water(time) ;
		neutral_wind_speed_relative_to_water:_FillValue = -9999. ;
		neutral_wind_speed_relative_to_water:long_name = "Neutral Wind Speed relative to water adjusted to 10m and neutral stratification computed from ADCP measurements" ;
		neutral_wind_speed_relative_to_water:valid_max = 13.3476314544678 ;
		neutral_wind_speed_relative_to_water:valid_min = 0. ;
		neutral_wind_speed_relative_to_water:add_offset = 0. ;
		neutral_wind_speed_relative_to_water:scale_factor = 1. ;
		neutral_wind_speed_relative_to_water:standard_name = "wind_speed" ;
		neutral_wind_speed_relative_to_water:units = "m s-1" ;
		neutral_wind_speed_relative_to_water:coverage_content_type = "physicalMeasurement" ;
		neutral_wind_speed_relative_to_water:coordinates = "time longitude latitude" ;
	double air_temperature_16p5m(time) ;
		air_temperature_16p5m:_FillValue = -9999. ;
		air_temperature_16p5m:long_name = "Air Temperature" ;
		air_temperature_16p5m:comment = "Air Temperature at ~16.5m from calibrated WHOI and UConn Air Temperature Sensors on the bow mast" ;
		air_temperature_16p5m:valid_max = 28.7145162081041 ;
		air_temperature_16p5m:valid_min = 23.1466122661809 ;
		air_temperature_16p5m:add_offset = 0. ;
		air_temperature_16p5m:scale_factor = 1. ;
		air_temperature_16p5m:standard_name = "air_temperature" ;
		air_temperature_16p5m:units = "degrees_C" ;
		air_temperature_16p5m:coverage_content_type = "physicalMeasurement" ;
		air_temperature_16p5m:coordinates = "time longitude latitude" ;
	double air_temperature(time) ;
		air_temperature:_FillValue = -9999. ;
		air_temperature:long_name = "Air Temperature" ;
		air_temperature:comment = "Air Temperature adjusted to 10m from calibrated WHOI and UConn Air Temperature Sensors on the bow mast" ;
		air_temperature:valid_max = 28.792594909668 ;
		air_temperature:valid_min = 23.2937183380127 ;
		air_temperature:add_offset = 0. ;
		air_temperature:scale_factor = 1. ;
		air_temperature:standard_name = "air_temperature" ;
		air_temperature:units = "degrees_C" ;
		air_temperature:coverage_content_type = "physicalMeasurement" ;
		air_temperature:coordinates = "time longitude latitude" ;
	double near_sea_surface_temperature_5cm(time) ;
		near_sea_surface_temperature_5cm:_FillValue = -9999. ;
		near_sea_surface_temperature_5cm:long_name = "Near Surface Sea Temperature at ~5cm from Sea-Snake after callibration with Osspre Sensors" ;
		near_sea_surface_temperature_5cm:valid_max = 32. ;
		near_sea_surface_temperature_5cm:valid_min = -1. ;
		near_sea_surface_temperature_5cm:add_offset = 0. ;
		near_sea_surface_temperature_5cm:scale_factor = 1. ;
		near_sea_surface_temperature_5cm:standard_name = "sea_water_temperature" ;
		near_sea_surface_temperature_5cm:units = "degrees_C" ;
		near_sea_surface_temperature_5cm:coverage_content_type = "physicalMeasurement" ;
		near_sea_surface_temperature_5cm:coordinates = "time longitude latitude" ;
	double near_sea_surface_temperature_2m(time) ;
		near_sea_surface_temperature_2m:_FillValue = -9999. ;
		near_sea_surface_temperature_2m:long_name = "Near Surface Sea Temperature at 2m from USPS" ;
		near_sea_surface_temperature_2m:valid_max = 32. ;
		near_sea_surface_temperature_2m:valid_min = -1. ;
		near_sea_surface_temperature_2m:add_offset = 0. ;
		near_sea_surface_temperature_2m:scale_factor = 1. ;
		near_sea_surface_temperature_2m:standard_name = "sea_water_temperature" ;
		near_sea_surface_temperature_2m:units = "degrees_C" ;
		near_sea_surface_temperature_2m:coverage_content_type = "physicalMeasurement" ;
		near_sea_surface_temperature_2m:coordinates = "time longitude latitude" ;
	double near_sea_surface_temperature_3m(time) ;
		near_sea_surface_temperature_3m:_FillValue = -9999. ;
		near_sea_surface_temperature_3m:long_name = "Near Surface Sea Temperature at 3m from USPS" ;
		near_sea_surface_temperature_3m:valid_max = 32. ;
		near_sea_surface_temperature_3m:valid_min = -1. ;
		near_sea_surface_temperature_3m:add_offset = 0. ;
		near_sea_surface_temperature_3m:scale_factor = 1. ;
		near_sea_surface_temperature_3m:standard_name = "sea_water_temperature" ;
		near_sea_surface_temperature_3m:units = "degrees_C" ;
		near_sea_surface_temperature_3m:coverage_content_type = "physicalMeasurement" ;
		near_sea_surface_temperature_3m:coordinates = "time longitude latitude" ;
	double near_sea_surface_temperature_5m(time) ;
		near_sea_surface_temperature_5m:_FillValue = -9999. ;
		near_sea_surface_temperature_5m:long_name = "Near Surface Sea Temperature at 5m from thermosalinograph" ;
		near_sea_surface_temperature_5m:valid_max = 32. ;
		near_sea_surface_temperature_5m:valid_min = -1. ;
		near_sea_surface_temperature_5m:add_offset = 0. ;
		near_sea_surface_temperature_5m:scale_factor = 1. ;
		near_sea_surface_temperature_5m:standard_name = "sea_water_temperature" ;
		near_sea_surface_temperature_5m:units = "degrees_C" ;
		near_sea_surface_temperature_5m:coverage_content_type = "physicalMeasurement" ;
		near_sea_surface_temperature_5m:coordinates = "time longitude latitude" ;
	double relative_humidity_16p5m(time) ;
		relative_humidity_16p5m:_FillValue = -9999. ;
		relative_humidity_16p5m:long_name = "Relative Humidity" ;
		relative_humidity_16p5m:comment = "Relative Humidity at ~16.5m reconstructed from Q, aspirated Tair, and P measurements" ;
		relative_humidity_16p5m:valid_max = 100. ;
		relative_humidity_16p5m:valid_min = 0. ;
		relative_humidity_16p5m:add_offset = 0. ;
		relative_humidity_16p5m:scale_factor = 1. ;
		relative_humidity_16p5m:standard_name = "relative_humidity" ;
		relative_humidity_16p5m:units = "%" ;
		relative_humidity_16p5m:coverage_content_type = "physicalMeasurement" ;
		relative_humidity_16p5m:coordinates = "time longitude latitude" ;
	double relative_humidity_2m(time) ;
		relative_humidity_2m:_FillValue = -9999. ;
		relative_humidity_2m:long_name = "Relative Humidity" ;
		relative_humidity_2m:comment = "Relative Humidity adjusted to 2m reconstructed from Q, aspirated Tair, and P measurements" ;
		relative_humidity_2m:valid_max = 100. ;
		relative_humidity_2m:valid_min = 0. ;
		relative_humidity_2m:add_offset = 0. ;
		relative_humidity_2m:scale_factor = 1. ;
		relative_humidity_2m:standard_name = "relative_humidity" ;
		relative_humidity_2m:units = "%" ;
		relative_humidity_2m:coverage_content_type = "physicalMeasurement" ;
		relative_humidity_2m:coordinates = "time longitude latitude" ;
	double relative_humidity_10m(time) ;
		relative_humidity_10m:_FillValue = -9999. ;
		relative_humidity_10m:long_name = "Relative Humidity" ;
		relative_humidity_10m:comment = "Relative Humidity adjusted to 10m reconstructed from Q, aspirated Tair, and P measurements" ;
		relative_humidity_10m:valid_max = 100. ;
		relative_humidity_10m:valid_min = 0. ;
		relative_humidity_10m:add_offset = 0. ;
		relative_humidity_10m:scale_factor = 1. ;
		relative_humidity_10m:standard_name = "relative_humidity" ;
		relative_humidity_10m:units = "%" ;
		relative_humidity_10m:coverage_content_type = "physicalMeasurement" ;
		relative_humidity_10m:coordinates = "time longitude latitude" ;
	double pressure(time) ;
		pressure:_FillValue = -9999. ;
		pressure:long_name = "Pressure from UConn Barometers on the 03 deck" ;
		pressure:valid_max = 1020. ;
		pressure:valid_min = 1000. ;
		pressure:add_offset = 0. ;
		pressure:scale_factor = 1. ;
		pressure:standard_name = "air_pressure" ;
		pressure:units = "mbar" ;
		pressure:coverage_content_type = "physicalMeasurement" ;
		pressure:coordinates = "time longitude latitude" ;
	double specific_humidity_16p5m(time) ;
		specific_humidity_16p5m:_FillValue = -9999. ;
		specific_humidity_16p5m:long_name = "Specific Humidity" ;
		specific_humidity_16p5m:comment = "Specific Humidity at ~16.5m computed from calibrated UConn and WHOI RH/T Sensors on the bow mast" ;
		specific_humidity_16p5m:valid_max = 20.4689352593528 ;
		specific_humidity_16p5m:valid_min = 13.0091783628398 ;
		specific_humidity_16p5m:add_offset = 0. ;
		specific_humidity_16p5m:scale_factor = 1. ;
		specific_humidity_16p5m:standard_name = "specific_humidity" ;
		specific_humidity_16p5m:units = "g kg-1" ;
		specific_humidity_16p5m:coverage_content_type = "physicalMeasurement" ;
		specific_humidity_16p5m:coordinates = "time longitude latitude" ;
	double specific_humidity_2m(time) ;
		specific_humidity_2m:_FillValue = -9999. ;
		specific_humidity_2m:long_name = "Specific Humidity" ;
		specific_humidity_2m:comment = "Specific Humidity adjusted to 2m computed from four Inter-Calibrated RH/T Sensors" ;
		specific_humidity_2m:valid_max = 20.8551940917969 ;
		specific_humidity_2m:valid_min = 14.242283821106 ;
		specific_humidity_2m:add_offset = 0. ;
		specific_humidity_2m:scale_factor = 1. ;
		specific_humidity_2m:standard_name = "specific_humidity" ;
		specific_humidity_2m:units = "g kg-1" ;
		specific_humidity_2m:coverage_content_type = "physicalMeasurement" ;
		specific_humidity_2m:coordinates = "time longitude latitude" ;
	double specific_humidity_10m(time) ;
		specific_humidity_10m:_FillValue = -9999. ;
		specific_humidity_10m:long_name = "Specific Humidity" ;
		specific_humidity_10m:comment = "Specific Humidity adjusted to 10m computed from four Inter-Calibrated RH/T Sensors" ;
		specific_humidity_10m:valid_max = 20.544979095459 ;
		specific_humidity_10m:valid_min = 13.2500047683716 ;
		specific_humidity_10m:add_offset = 0. ;
		specific_humidity_10m:scale_factor = 1. ;
		specific_humidity_10m:standard_name = "specific_humidity" ;
		specific_humidity_10m:units = "g kg-1" ;
		specific_humidity_10m:coverage_content_type = "physicalMeasurement" ;
		specific_humidity_10m:coordinates = "time longitude latitude" ;
	double specific_humidity_sea_surface(time) ;
		specific_humidity_sea_surface:_FillValue = -9999. ;
		specific_humidity_sea_surface:long_name = "Specific Humidity at Sea Surface" ;
		specific_humidity_sea_surface:comment = "Specific Humidity at Sea Surface computed from SST" ;
		specific_humidity_sea_surface:valid_max = 28.1663436889648 ;
		specific_humidity_sea_surface:valid_min = 21.5090866088867 ;
		specific_humidity_sea_surface:add_offset = 0. ;
		specific_humidity_sea_surface:scale_factor = 1. ;
		specific_humidity_sea_surface:standard_name = "surface_specific_humidity" ;
		specific_humidity_sea_surface:units = "g kg-1" ;
		specific_humidity_sea_surface:coverage_content_type = "physicalMeasurement" ;
		specific_humidity_sea_surface:coordinates = "time longitude latitude" ;
	double sss(time) ;
		sss:_FillValue = -9999. ;
		sss:long_name = "Sea surface salinity from the salinity snake" ;
		sss:valid_max = 42. ;
		sss:valid_min = 2. ;
		sss:add_offset = 0. ;
		sss:scale_factor = 1. ;
		sss:standard_name = "sea_surface_salinity" ;
		sss:units = "1" ;
		sss:coverage_content_type = "physicalMeasurement" ;
		sss:coordinates = "time longitude latitude" ;
	double salinity_2m(time) ;
		salinity_2m:_FillValue = -9999. ;
		salinity_2m:long_name = "Salinity at 2m from USPS" ;
		salinity_2m:valid_max = 42. ;
		salinity_2m:valid_min = 2. ;
		salinity_2m:add_offset = 0. ;
		salinity_2m:scale_factor = 1. ;
		salinity_2m:standard_name = "sea_water_practical_salinity" ;
		salinity_2m:units = "1" ;
		salinity_2m:coverage_content_type = "physicalMeasurement" ;
		salinity_2m:coordinates = "time longitude latitude" ;
	double salinity_3m(time) ;
		salinity_3m:_FillValue = -9999. ;
		salinity_3m:long_name = "Salinity at 3m from USPS" ;
		salinity_3m:valid_max = 42. ;
		salinity_3m:valid_min = 2. ;
		salinity_3m:add_offset = 0. ;
		salinity_3m:scale_factor = 1. ;
		salinity_3m:standard_name = "sea_water_practical_salinity" ;
		salinity_3m:units = "1" ;
		salinity_3m:coverage_content_type = "physicalMeasurement" ;
		salinity_3m:coordinates = "time longitude latitude" ;
	double salinity_5m(time) ;
		salinity_5m:_FillValue = -9999. ;
		salinity_5m:long_name = "Salinity at 5m from thermosalinograph" ;
		salinity_5m:valid_max = 42. ;
		salinity_5m:valid_min = 2. ;
		salinity_5m:add_offset = 0. ;
		salinity_5m:scale_factor = 1. ;
		salinity_5m:standard_name = "sea_water_practical_salinity" ;
		salinity_5m:units = "1" ;
		salinity_5m:coverage_content_type = "physicalMeasurement" ;
		salinity_5m:coordinates = "time longitude latitude" ;
	double precipitation_rate(time) ;
		precipitation_rate:_FillValue = -9999. ;
		precipitation_rate:long_name = "Precipitation rate of Optical Rain Gauge" ;
		precipitation_rate:valid_max = 150. ;
		precipitation_rate:valid_min = 0. ;
		precipitation_rate:add_offset = 0. ;
		precipitation_rate:scale_factor = 1. ;
		precipitation_rate:standard_name = "lwe_precipitation_rate" ;
		precipitation_rate:units = "mm hr-1" ;
		precipitation_rate:coverage_content_type = "physicalMeasurement" ;
		precipitation_rate:coordinates = "time longitude latitude" ;
	double evaporation_rate(time) ;
		evaporation_rate:_FillValue = -9999. ;
		evaporation_rate:long_name = "Evaporation rate of Optical Rain Gauge" ;
		evaporation_rate:valid_max = 2. ;
		evaporation_rate:valid_min = 0. ;
		evaporation_rate:add_offset = 0. ;
		evaporation_rate:scale_factor = 1. ;
		evaporation_rate:standard_name = "lwe_water_evaporation_rate" ;
		evaporation_rate:units = "mm hr-1" ;
		evaporation_rate:coverage_content_type = "physicalMeasurement" ;
		evaporation_rate:coordinates = "time longitude latitude" ;

// global attributes:
		:DOI = "10.5067/SMODE-RVMET" ;
		:title = "S-MODE Pilot Field Campaign Fall 2020 Shipboard Meteorology measurements from the R/V Oceanus<, XXXX>" ;
		:summary = "S-MODE Pilot Field Campaign Fall 2020 Shipboard Meteorology measurements from the R/V Oceanus<, XXXX>" ;
		:keywords = "EARTH SCIENCE > OCEANS > SALINITY/DENSITY > CONDUCTIVITY, EARTH SCIENCE > OCEANS > PRECIPITATION > PRECIPITATION RATE, EARTH SCIENCE > OCEANS > OCEAN WINDS > SURFACE WINDS > WIND DIRECTION, EARTH SCIENCE > OCEANS > OCEAN WINDS > SURFACE WINDS > WIND SPEED, EARTH SCIENCE > OCEANS > SALINITY/DENSITY > SALINITY, EARTH SCIENCE > OCEANS > OCEAN TEMPERATURE > SEA SURFACE TEMPERATURE, EARTH SCIENCE > ATMOSPHERE > ATMOSPHERIC PRESSURE > ATMOSPHERIC PRESSURE MEASUREMENTS, EARTH SCIENCE > ATMOSPHERE > ATMOSPHERIC TEMPERATURE > SURFACE TEMPERATURE" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:conventions = "CF-1.8, ACDD-1.3" ;
		:id = "PODAAC-SMODE-RVMET" ;
		:uuid = "7d5a12d7-17b3-460c-be43-1ec2af2a33b2" ;
		:naming_authority = "gov.nasa" ;
		:featureType = "trajectory" ;
		:cdm_data_type = "Trajectory" ;
		:source = "S-MODE_PFC_OC2004B_meteorology_##.nc.cdl" ;
		:platform = "In Situ Ocean-based Platforms > SHIPS > RV Oceanus" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:instrument = "In Situ/Laboratory Instruments > Recorders/Loggers > > > MMS" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:processing_level = "L2" ;
		:standard_name_vocabulary = "CF Standard Name Table v72" ;
		:acknowledgement = "TBD" ;
		:comment = "" ;
		:license = "S-MODE data are considered experimental and not to be used for any purpose for which life or property is potentially at risk. Distributor assumes no responsibility for the manner in which the data are used. Otherwise data are free for public use." ;
		:product_version = "1" ;
		:metadata_link = "https://doi.org/10.5067/SMODE-RVMET" ;
		:creator_name = "Melissa Omand" ;
		:creator_email = "momand@uri.edu" ;
		:creator_type = "person" ;
		:creator_institution = "URI/" ;
		:institution = "URI/" ;
		:project = "Sub-Mesoscale Ocean Dynamics Experiment (S-MODE)" ;
		:program = "NASA Earth Venture Suborbital-3 (EVS-3)" ;
		:contributor_name = "Frederick Bingham" ;
		:contributor_role = "Project Data Manager" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center, Jet Propulsion Laboratory, NASA" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:sea_name = "Pacific" ;
		:geospatial_lat_min = 5.06140075 ;
		:geospatial_lat_max = 13.4568725 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = "0.1 degrees" ;
		:geospatial_lon_min = -144.87482775 ;
		:geospatial_lon_max = -123.37702175 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = "0.1 degrees" ;
		:geospatial_vertical_min = 1006.588 ;
		:geospatial_vertical_max = 1014.882 ;
		:geospatial_vertical_resolution = "1 meters" ;
		:geospatial_vertical_units = "meters" ;
		:geospatial_vertical_positive = "down" ;
		:time_coverage_start = "2016-08-20T00:00:30" ;
		:time_coverage_end = "2016-09-18T23:59:30" ;
		:date_created = "2020-09-01T14:11:36" ;
}
