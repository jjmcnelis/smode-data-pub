netcdf prm20160125t195943_refl {
dimensions:
	x = 197 ;
	y = 985 ;
	band = 246 ;
variables:
	double x(x) ;
		x:units = "m" ;
		x:axis = "X" ;
		x:standard_name = "projection_x_coordinate" ;
		x:long_name = "x coordinate of projection" ;
	double y(y) ;
		y:units = "m" ;
		y:axis = "Y" ;
		y:standard_name = "projection_y_coordinate" ;
		y:long_name = "y coordinate of projection" ;
	float lat(y, x) ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
	float lon(y, x) ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
	char UTM_Projection ;
		UTM_Projection:crs_wkt = "PROJCRS[\"unknown\",BASEGEOGCRS[\"unknown\",DATUM[\"World Geodetic System 1984\",ELLIPSOID[\"WGS 84\",6378137,298.257223563,LENGTHUNIT[\"metre\",1]],ID[\"EPSG\",6326]],PRIMEM[\"Greenwich\",0,ANGLEUNIT[\"degree\",0.0174532925199433],ID[\"EPSG\",8901]]],CONVERSION[\"UTM zone 19S\",METHOD[\"Transverse Mercator\",ID[\"EPSG\",9807]],PARAMETER[\"Latitude of natural origin\",0,ANGLEUNIT[\"degree\",0.0174532925199433],ID[\"EPSG\",8801]],PARAMETER[\"Longitude of natural origin\",-69,ANGLEUNIT[\"degree\",0.0174532925199433],ID[\"EPSG\",8802]],PARAMETER[\"Scale factor at natural origin\",0.9996,SCALEUNIT[\"unity\",1],ID[\"EPSG\",8805]],PARAMETER[\"False easting\",500000,LENGTHUNIT[\"metre\",1],ID[\"EPSG\",8806]],PARAMETER[\"False northing\",10000000,LENGTHUNIT[\"metre\",1],ID[\"EPSG\",8807]],ID[\"EPSG\",17019]],CS[Cartesian,2],AXIS[\"(E)\",east,ORDER[1],LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]]],AXIS[\"(N)\",north,ORDER[2],LENGTHUNIT[\"metre\",1,ID[\"EPSG\",9001]]]]" ;
		UTM_Projection:semi_major_axis = 6378137. ;
		UTM_Projection:semi_minor_axis = 6356752.31424518 ;
		UTM_Projection:inverse_flattening = 298.257223563 ;
		UTM_Projection:reference_ellipsoid_name = "WGS 84" ;
		UTM_Projection:longitude_of_prime_meridian = 0. ;
		UTM_Projection:prime_meridian_name = "Greenwich" ;
		UTM_Projection:geographic_crs_name = "unknown" ;
		UTM_Projection:horizontal_datum_name = "World Geodetic System 1984" ;
		UTM_Projection:projected_crs_name = "unknown" ;
		UTM_Projection:grid_mapping_name = "transverse_mercator" ;
		UTM_Projection:latitude_of_projection_origin = 0. ;
		UTM_Projection:longitude_of_central_meridian = -69. ;
		UTM_Projection:false_easting = 500000. ;
		UTM_Projection:false_northing = 10000000. ;
		UTM_Projection:scale_factor_at_central_meridian = 0.9996 ;
	float wavelength(band) ;
		wavelength:long_name = "wavelengths of band centers" ;
		wavelength:units = "nm" ;
		wavelength:valid_min = 350.f ;
		wavelength:valid_max = 1050.f ;
	float correction_factors(band) ;
		correction_factors:long_name = "correction factors" ;
		correction_factors:units = "unitless" ;
		correction_factors:valid_min = 1.f ;
		correction_factors:valid_max = 1.f ;
	float reflectance(band, y, x) ;
		reflectance:_FillValue = -9999.f ;
		reflectance:long_name = "reflectance" ;
		reflectance:units = "unitless" ;
		reflectance:valid_min = 0. ;
		reflectance:valid_max = 1000. ;
		reflectance:grid_mapping = "UTM_Projection" ;
		reflectance:coordinates = "lat lon" ;

// global attributes:
		:id = "10.5067/PRISM/#" ;
		:naming_authority = "gov.nasa.jpl.prism" ;
		:license = "https://science.nasa.gov/earth-science/earth-science-data/data-information-policy/" ;
		:project = "NASA PRISM" ;
		:project_url = "https://prism.jpl.nasa.gov/" ;
		:institution = "NASA Jet Propulsion Laboratory" ;
		:instrument = "PRISM (Portable Remote Imaging SpectroMeter)" ;
		:platform = "G-IV (Gulfstream-IV)" ;
		:Conventions = "CF-1.7" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:standard_name_vocabulary = "CF Standard Names v72" ;
		:processing_version = "V1.0" ;
		:product_version = "v1w2" ;
		:product_name = "prm20160125t195943_refl.nc" ;
		:creator_name = "PRISM Science Team" ;
		:creator_role = "group" ;
		:creator_url = "https://prism.jpl.nasa.gov" ;
		:creator_email = "sarah.r.lundeen@jpl.nasa.gov" ;
		:publisher_name = "PRISM Science Team" ;
		:publisher_role = "group" ;
		:publisher_url = "https://prism.jpl.nasa.gov" ;
		:publisher_email = "sarah.r.lundeen@jpl.nasa.gov" ;
		:date_created = "2020-08-25T08:46:36Z" ;
		:date_updated = "2020-08-25T08:46:36Z" ;
		:geospatial_lon_min = -69.5124713973911 ;
		:geospatial_lon_max = -69.4649447642403 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lat_min = -67.8077637789882 ;
		:geospatial_lat_max = -67.7206939671764 ;
		:geospatial_lat_units = "degrees_north" ;
		:title = "PRISM Level-2 Reflectance" ;
		:processing_level = "L2" ;
}
