netcdf S-MODE_PFC_OC2004B_thermosalinograph_\#\# {
dimensions:
	time = 673920 ;
variables:
	double time(time) ;
		time:long_name = "Time of Underway Salinity Profiling System measurement" ;
		time:axis = "T" ;
		time:standard_name = "time" ;
		time:units = "days since 1950-01-01 00:00:00" ;
		time:coverage_content_type = "coordinate" ;
	double longitude(time) ;
		longitude:_FillValue = -9999. ;
		longitude:long_name = "Longitude of Underway Salinity Profiling System measurement" ;
		longitude:valid_max = 180. ;
		longitude:valid_min = -180. ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "referenceInformation" ;
	double latitude(time) ;
		latitude:_FillValue = -9999. ;
		latitude:long_name = "Latitude of Underway Salinity Profiling System measurement" ;
		latitude:valid_max = 90. ;
		latitude:valid_min = -90. ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "referenceInformation" ;
	double speed_over_ground(time) ;
		speed_over_ground:_FillValue = -9999. ;
		speed_over_ground:long_name = "Speed Over Ground of Underway Salinity Profiling System measurement" ;
		speed_over_ground:valid_max = 20. ;
		speed_over_ground:valid_min = 0. ;
		speed_over_ground:add_offset = 0. ;
		speed_over_ground:scale_factor = 1. ;
		speed_over_ground:standard_name = "platform_speed_wrt_ground" ;
		speed_over_ground:units = "m s-1" ;
		speed_over_ground:coverage_content_type = "physicalMeasurement" ;
		speed_over_ground:coordinates = "time longitude latitude" ;
	double course_over_ground(time) ;
		course_over_ground:_FillValue = -9999. ;
		course_over_ground:long_name = "Course Over Ground of Underway Salinity Profiling System measurement" ;
		course_over_ground:valid_max = 360. ;
		course_over_ground:valid_min = 0. ;
		course_over_ground:add_offset = 0. ;
		course_over_ground:scale_factor = 1. ;
		course_over_ground:standard_name = "platform_course" ;
		course_over_ground:units = "degrees" ;
		course_over_ground:coverage_content_type = "physicalMeasurement" ;
		course_over_ground:coordinates = "time longitude latitude" ;
	double pressure_2m(time) ;
		pressure_2m:_FillValue = -9999. ;
		pressure_2m:long_name = "Pressure at 2m of Underway Salinity Profiling System measurement" ;
		pressure_2m:valid_max = 10. ;
		pressure_2m:valid_min = 0. ;
		pressure_2m:add_offset = 0. ;
		pressure_2m:scale_factor = 1. ;
		pressure_2m:standard_name = "sea_water_pressure" ;
		pressure_2m:units = "dbar" ;
		pressure_2m:coverage_content_type = "physicalMeasurement" ;
		pressure_2m:coordinates = "time longitude latitude" ;
	double pressure_3m(time) ;
		pressure_3m:_FillValue = -9999. ;
		pressure_3m:long_name = "Pressure at 3m of Underway Salinity Profiling System measurement" ;
		pressure_3m:valid_max = 10. ;
		pressure_3m:valid_min = 0. ;
		pressure_3m:add_offset = 0. ;
		pressure_3m:scale_factor = 1. ;
		pressure_3m:standard_name = "sea_water_pressure" ;
		pressure_3m:units = "dbar" ;
		pressure_3m:coverage_content_type = "physicalMeasurement" ;
		pressure_3m:coordinates = "time longitude latitude" ;
	double density_2m(time) ;
		density_2m:_FillValue = -9999. ;
		density_2m:long_name = "Density at 2m of Underway Salinity Profiling System measurement" ;
		density_2m:valid_max = 1030. ;
		density_2m:valid_min = 1010. ;
		density_2m:add_offset = 0. ;
		density_2m:coordinates = "time longitude latitude" ;
		density_2m:scale_factor = 1. ;
		density_2m:standard_name = "sea_water_density" ;
		density_2m:units = "kg m-3" ;
		density_2m:coverage_content_type = "physicalMeasurement" ;
	double density_3m(time) ;
		density_3m:_FillValue = -9999. ;
		density_3m:long_name = "Density at 3m of Underway Salinity Profiling System measurement" ;
		density_3m:valid_max = 1030. ;
		density_3m:valid_min = 1010. ;
		density_3m:add_offset = 0. ;
		density_3m:coordinates = "time longitude latitude" ;
		density_3m:scale_factor = 1. ;
		density_3m:standard_name = "sea_water_density" ;
		density_3m:units = "kg m-3" ;
		density_3m:coverage_content_type = "physicalMeasurement" ;
	double salinity_2m(time) ;
		salinity_2m:_FillValue = -9999. ;
		salinity_2m:long_name = "Salinity at 2m of Underway Salinity Profiling System measurement" ;
		salinity_2m:valid_max = 42. ;
		salinity_2m:valid_min = 2. ;
		salinity_2m:add_offset = 0. ;
		salinity_2m:scale_factor = 1. ;
		salinity_2m:standard_name = "sea_water_practical_salinity" ;
		salinity_2m:units = "1" ;
		salinity_2m:coverage_content_type = "physicalMeasurement" ;
		salinity_2m:coordinates = "time longitude latitude" ;
	double salinity_3m(time) ;
		salinity_3m:_FillValue = -9999. ;
		salinity_3m:long_name = "Salinity at 3m of Underway Salinity Profiling System measurement" ;
		salinity_3m:valid_max = 42. ;
		salinity_3m:valid_min = 2. ;
		salinity_3m:add_offset = 0. ;
		salinity_3m:scale_factor = 1. ;
		salinity_3m:standard_name = "sea_water_practical_salinity" ;
		salinity_3m:units = "1" ;
		salinity_3m:coverage_content_type = "physicalMeasurement" ;
		salinity_3m:coordinates = "time longitude latitude" ;
	double uncorrected_salinity_5m(time) ;
		uncorrected_salinity_5m:_FillValue = -9999. ;
		uncorrected_salinity_5m:long_name = "Uncorrected Salinity at 5m of Underway Salinity Profiling System measurement" ;
		uncorrected_salinity_5m:valid_max = 42. ;
		uncorrected_salinity_5m:valid_min = 2. ;
		uncorrected_salinity_5m:add_offset = 0. ;
		uncorrected_salinity_5m:scale_factor = 1. ;
		uncorrected_salinity_5m:standard_name = "sea_water_practical_salinity" ;
		uncorrected_salinity_5m:units = "1" ;
		uncorrected_salinity_5m:coverage_content_type = "physicalMeasurement" ;
		uncorrected_salinity_5m:coordinates = "time longitude latitude" ;
	double temperature_2m(time) ;
		temperature_2m:_FillValue = -9999. ;
		temperature_2m:long_name = "Temperature at 2m of Underway Salinity Profiling System measurement" ;
		temperature_2m:valid_max = 32. ;
		temperature_2m:valid_min = -1. ;
		temperature_2m:add_offset = 0. ;
		temperature_2m:scale_factor = 1. ;
		temperature_2m:standard_name = "sea_water_temperature" ;
		temperature_2m:units = "degrees_C" ;
		temperature_2m:coverage_content_type = "physicalMeasurement" ;
		temperature_2m:coordinates = "time longitude latitude" ;
	double temperature_3m(time) ;
		temperature_3m:_FillValue = -9999. ;
		temperature_3m:long_name = "Temperature at 3m of Underway Salinity Profiling System measurement" ;
		temperature_3m:valid_max = 32. ;
		temperature_3m:valid_min = -1. ;
		temperature_3m:add_offset = 0. ;
		temperature_3m:scale_factor = 1. ;
		temperature_3m:standard_name = "sea_water_temperature" ;
		temperature_3m:units = "degrees_C" ;
		temperature_3m:coverage_content_type = "physicalMeasurement" ;
		temperature_3m:coordinates = "time longitude latitude" ;
	double uncorrected_temperature_5m(time) ;
		uncorrected_temperature_5m:_FillValue = -9999. ;
		uncorrected_temperature_5m:long_name = "Uncorrected Temperature at 5m of Underway Salinity Profiling System measurement" ;
		uncorrected_temperature_5m:valid_max = 32. ;
		uncorrected_temperature_5m:valid_min = -1. ;
		uncorrected_temperature_5m:add_offset = 0. ;
		uncorrected_temperature_5m:scale_factor = 1. ;
		uncorrected_temperature_5m:standard_name = "sea_water_temperature" ;
		uncorrected_temperature_5m:units = "degrees_C" ;
		uncorrected_temperature_5m:coverage_content_type = "physicalMeasurement" ;
		uncorrected_temperature_5m:coordinates = "time longitude latitude" ;
	double downwelling_longwave_infrared_radiation(time) ;
		downwelling_longwave_infrared_radiation:_FillValue = -9999. ;
		downwelling_longwave_infrared_radiation:long_name = "Downwelling Longwave (infrared) Radiation" ;
		downwelling_longwave_infrared_radiation:valid_max = 600. ;
		downwelling_longwave_infrared_radiation:valid_min = 0. ;
		downwelling_longwave_infrared_radiation:add_offset = 0. ;
		downwelling_longwave_infrared_radiation:scale_factor = 1. ;
		downwelling_longwave_infrared_radiation:standard_name = "downwelling_longwave_radiance_in_air" ;
		downwelling_longwave_infrared_radiation:units = "W m-2" ;
		downwelling_longwave_infrared_radiation:coverage_content_type = "physicalMeasurement" ;
		downwelling_longwave_infrared_radiation:coordinates = "time longitude latitude" ;
	double downwelling_shortwave_solar_radiation(time) ;
		downwelling_shortwave_solar_radiation:_FillValue = -9999. ;
		downwelling_shortwave_solar_radiation:long_name = "Downwelling Shortwave (solar) Radiation" ;
		downwelling_shortwave_solar_radiation:valid_max = 1500. ;
		downwelling_shortwave_solar_radiation:valid_min = 0. ;
		downwelling_shortwave_solar_radiation:add_offset = 0. ;
		downwelling_shortwave_solar_radiation:scale_factor = 1. ;
		downwelling_shortwave_solar_radiation:standard_name = "downwelling_shortwave_radiance_in_air" ;
		downwelling_shortwave_solar_radiation:units = "W m-2" ;
		downwelling_shortwave_solar_radiation:coverage_content_type = "physicalMeasurement" ;
		downwelling_shortwave_solar_radiation:coordinates = "time longitude latitude" ;
	double relative_humidity(time) ;
		relative_humidity:_FillValue = -9999. ;
		relative_humidity:long_name = "Relative Humidity" ;
		relative_humidity:valid_max = 100. ;
		relative_humidity:valid_min = 0. ;
		relative_humidity:add_offset = 0. ;
		relative_humidity:scale_factor = 1. ;
		relative_humidity:standard_name = "relative_humidity" ;
		relative_humidity:units = "%" ;
		relative_humidity:coverage_content_type = "physicalMeasurement" ;
		relative_humidity:coordinates = "time longitude latitude" ;
	double cumulative_rain(time) ;
		cumulative_rain:_FillValue = -9999. ;
		cumulative_rain:long_name = "Cumulative Rain" ;
		cumulative_rain:valid_max = 100. ;
		cumulative_rain:valid_min = 0. ;
		cumulative_rain:add_offset = 0. ;
		cumulative_rain:scale_factor = 1. ;
		cumulative_rain:standard_name = "thickness_of_rainfall_amount" ;
		cumulative_rain:units = "mm" ;
		cumulative_rain:coverage_content_type = "physicalMeasurement" ;
		cumulative_rain:coordinates = "time longitude latitude" ;
	double wind_direction(time) ;
		wind_direction:_FillValue = -9999. ;
		wind_direction:long_name = "True Wind Direction at about 17 m above sea level (direction wind came from)" ;
		wind_direction:valid_max = 360. ;
		wind_direction:valid_min = 0. ;
		wind_direction:add_offset = 0. ;
		wind_direction:scale_factor = 1. ;
		wind_direction:standard_name = "wind_from_direction" ;
		wind_direction:units = "degree" ;
		wind_direction:coverage_content_type = "physicalMeasurement" ;
		wind_direction:coordinates = "time longitude latitude" ;
	double wind_speed(time) ;
		wind_speed:_FillValue = -9999. ;
		wind_speed:long_name = "Wind Speed" ;
		wind_speed:valid_max = 50. ;
		wind_speed:valid_min = 0. ;
		wind_speed:add_offset = 0. ;
		wind_speed:scale_factor = 1. ;
		wind_speed:standard_name = "wind_speed" ;
		wind_speed:units = "m s-1" ;
		wind_speed:coverage_content_type = "physicalMeasurement" ;
		wind_speed:coordinates = "time longitude latitude" ;
	double ship_heave(time) ;
		ship_heave:_FillValue = -9999. ;
		ship_heave:long_name = "Ship Heave" ;
		ship_heave:valid_max = 1.96 ;
		ship_heave:valid_min = -1.82533270122604 ;
		ship_heave:add_offset = 0. ;
		ship_heave:scale_factor = 1. ;
		ship_heave:standard_name = "platform_heave" ;
		ship_heave:units = "m" ;
		ship_heave:coverage_content_type = "physicalMeasurement" ;
		ship_heave:coordinates = "time longitude latitude" ;
	double ship_pitch(time) ;
		ship_pitch:_FillValue = -9999. ;
		ship_pitch:long_name = "Ship Pitch Angle" ;
		ship_pitch:valid_max = 3.93533491404861 ;
		ship_pitch:valid_min = -3.92866468898443 ;
		ship_pitch:add_offset = 0. ;
		ship_pitch:scale_factor = 1. ;
		ship_pitch:standard_name = "platform_pitch_angle" ;
		ship_pitch:units = "degree" ;
		ship_pitch:coverage_content_type = "physicalMeasurement" ;
		ship_pitch:coordinates = "time longitude latitude" ;
	double ship_roll(time) ;
		ship_roll:_FillValue = -9999. ;
		ship_roll:long_name = "Ship Roll Angle" ;
		ship_roll:valid_max = 5.58933365877471 ;
		ship_roll:valid_min = -6.68800035941603 ;
		ship_roll:add_offset = 0. ;
		ship_roll:scale_factor = 1. ;
		ship_roll:standard_name = "platform_roll_angle" ;
		ship_roll:units = "degree" ;
		ship_roll:coverage_content_type = "physicalMeasurement" ;
		ship_roll:coordinates = "time longitude latitude" ;
	double air_pressure(time) ;
		air_pressure:_FillValue = -9999. ;
		air_pressure:long_name = "Air Pressure" ;
		air_pressure:valid_max = 1020. ;
		air_pressure:valid_min = 1000. ;
		air_pressure:add_offset = 0. ;
		air_pressure:scale_factor = 1. ;
		air_pressure:standard_name = "air_pressure" ;
		air_pressure:units = "mbar" ;
		air_pressure:coverage_content_type = "physicalMeasurement" ;
		air_pressure:coordinates = "time longitude latitude" ;
	double air_temperature(time) ;
		air_temperature:_FillValue = -9999. ;
		air_temperature:long_name = "Air Temperature" ;
		air_temperature:valid_max = 40. ;
		air_temperature:valid_min = 0. ;
		air_temperature:add_offset = 0. ;
		air_temperature:scale_factor = 1. ;
		air_temperature:standard_name = "air_temperature" ;
		air_temperature:units = "degrees_C" ;
		air_temperature:coverage_content_type = "physicalMeasurement" ;
		air_temperature:coordinates = "time longitude latitude" ;

// global attributes:
		:DOI = "10.5067/SMODE-RVTSG" ;
		:title = "S-MODE Pilot Field Campaign Fall 2020 Shipboard Thermosalinograph Measurements from R/V Oceanus<, XXXX>" ;
		:summary = "S-MODE Pilot Field Campaign Fall 2020 Shipboard Thermosalinograph Measurements from R/V Oceanus<, XXXX>" ;
		:keywords = "EARTH SCIENCE > OCEANS > SALINITY/DENSITY > CONDUCTIVITY, EARTH SCIENCE > OCEANS > PRECIPITATION > PRECIPITATION RATE, EARTH SCIENCE > OCEANS > OCEAN WINDS > SURFACE WINDS > WIND SPEED, EARTH SCIENCE > OCEANS > OCEAN WINDS > SURFACE WINDS > WIND DIRECTION, EARTH SCIENCE > OCEANS > SALINITY/DENSITY > SALINITY, EARTH SCIENCE > OCEANS > OCEAN TEMPERATURE > SEA SURFACE TEMPERATURE" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:conventions = "CF-1.8, ACDD-1.3" ;
		:id = "PODAAC-SMODE-RVTSG" ;
		:uuid = "ccdf6e87-f99a-4907-a4b4-56fcc6be8ab2" ;
		:naming_authority = "gov.nasa" ;
		:featureType = "trajectory" ;
		:cdm_data_type = "Trajectory" ;
		:source = "S-MODE_PFC_OC2004B_thermosalinograph_##.nc.cdl" ;
		:platform = "In Situ Ocean-based Platforms > SHIPS > RV Oceanus" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:instrument = "In Situ/Laboratory Instruments > Profilers/Sounders > > > THERMOSALINOGRAPHS" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:processing_level = "L2" ;
		:standard_name_vocabulary = "CF Standard Name Table v72" ;
		:acknowledgement = "TBD" ;
		:comment = "" ;
		:license = "S-MODE data are considered experimental and not to be used for any purpose for which life or property is potentially at risk. Distributor assumes no responsibility for the manner in which the data are used. Otherwise data are free for public use." ;
		:product_version = "1" ;
		:metadata_link = "https://doi.org/10.5067/SMODE-RVTSG" ;
		:creator_name = "Melissa Omand" ;
		:creator_email = "momand@uri.edu" ;
		:creator_type = "person" ;
		:creator_institution = "URI/" ;
		:institution = "URI/" ;
		:project = "Sub-Mesoscale Ocean Dynamics Experiment (S-MODE)" ;
		:program = "NASA Earth Venture Suborbital-3 (EVS-3)" ;
		:contributor_name = "Frederick Bingham" ;
		:contributor_role = "Project Data Manager" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center, Jet Propulsion Laboratory, NASA" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:sea_name = "Pacific" ;
		:geospatial_lat_min = 5.061344 ;
		:geospatial_lat_max = 18.6293995333687 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = "0.1 degrees" ;
		:geospatial_lon_min = -157.110813733344 ;
		:geospatial_lon_max = -123.377014266668 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = "0.1 degrees" ;
		:geospatial_vertical_min = 2. ;
		:geospatial_vertical_max = 5. ;
		:geospatial_vertical_resolution = "1 meters" ;
		:geospatial_vertical_units = "meters" ;
		:geospatial_vertical_positive = "down" ;
		:time_coverage_start = "YYYY-MM-DDTHH:MM:SS" ;
		:time_coverage_end = "2016-09-22T23:59:55" ;
		:date_created = "2020-09-01T14:19:07" ;
}
