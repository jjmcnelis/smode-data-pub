3,4c3,4
< 	time = 1 ;
< 	depth = 79246 ;
---
> 	time = 79246 ;
> 	timeSeries = 1 ;
5a6,8
>     int platform_id(timeSeries) ;
>         platform_id:long_name = "Unique identifier for each platform's time series  " ;
>         platform_id:cf_role = "timeseries_id" ;
12,13c15
< 	double latitude(time) ;
< 		latitude:_FillValue = NaN ;
---
> 	double latitude(timeSeries) ;
15,17d16
< 		latitude:valid_max = 90. ;
< 		latitude:valid_min = -90. ;
< 		latitude:axis = "Y" ;
20,22c19,20
< 		latitude:coverage_content_type = "coordinate" ;
< 	double longitude(time) ;
< 		longitude:_FillValue = NaN ;
---
> 		latitude:coverage_content_type = "referenceInformation" ;
> 	double longitude(timeSeries) ;
24,26d21
< 		longitude:valid_max = 180. ;
< 		longitude:valid_min = -180. ;
< 		longitude:axis = "X" ;
29,31c24,25
< 		longitude:coverage_content_type = "coordinate" ;
< 	double depth(depth) ;
< 		depth:_FillValue = NaN ;
---
> 		longitude:coverage_content_type = "referenceInformation" ;
> 	double depth(time) ;
35d28
< 		depth:axis = "Z" ;
39,224c32,205
< 		depth:coverage_content_type = "coordinate" ;
< 	double pressure(depth) ;
< 		pressure:_FillValue = NaN ;
< 		pressure:long_name = "Pressure of CTD measurement" ;
< 		pressure:valid_max = 1500. ;
< 		pressure:valid_min = -1. ;
< 		pressure:add_offset = 0. ;
< 		pressure:coordinates = "time depth latitude longitude" ;
< 		pressure:scale_factor = 1. ;
< 		pressure:standard_name = "sea_water_pressure" ;
< 		pressure:units = "dbar" ;
< 		pressure:coverage_content_type = "physicalMeasurement" ;
< 	double temperature(depth) ;
< 		temperature:_FillValue = NaN ;
< 		temperature:long_name = "Temperature of CTD measurement" ;
< 		temperature:valid_max = 32. ;
< 		temperature:valid_min = -1. ;
< 		temperature:add_offset = 0. ;
< 		temperature:coordinates = "time depth latitude longitude" ;
< 		temperature:scale_factor = 1. ;
< 		temperature:standard_name = "sea_water_temperature" ;
< 		temperature:units = "degrees_C" ;
< 		temperature:coverage_content_type = "physicalMeasurement" ;
< 	double temperature2(depth) ;
< 		temperature2:_FillValue = NaN ;
< 		temperature2:long_name = "Temperature of second CTD measurement" ;
< 		temperature2:valid_max = 32. ;
< 		temperature2:valid_min = -1. ;
< 		temperature2:add_offset = 0. ;
< 		temperature2:coordinates = "time depth latitude longitude" ;
< 		temperature2:scale_factor = 1. ;
< 		temperature2:standard_name = "sea_water_temperature" ;
< 		temperature2:units = "degrees_C" ;
< 		temperature2:coverage_content_type = "physicalMeasurement" ;
< 	double conductivity(depth) ;
< 		conductivity:_FillValue = NaN ;
< 		conductivity:long_name = "Conductivity of CTD measurement" ;
< 		conductivity:valid_max = 60. ;
< 		conductivity:valid_min = 0. ;
< 		conductivity:add_offset = 0. ;
< 		conductivity:coordinates = "time depth latitude longitude" ;
< 		conductivity:scale_factor = 1. ;
< 		conductivity:standard_name = "sea_water_electrical_conductivity" ;
< 		conductivity:units = "S m-1" ;
< 		conductivity:coverage_content_type = "physicalMeasurement" ;
< 	double conductivity2(depth) ;
< 		conductivity2:_FillValue = NaN ;
< 		conductivity2:long_name = "Conductivity of second CTD measurement" ;
< 		conductivity2:valid_max = 60. ;
< 		conductivity2:valid_min = 0. ;
< 		conductivity2:add_offset = 0. ;
< 		conductivity2:coordinates = "time depth latitude longitude" ;
< 		conductivity2:scale_factor = 1. ;
< 		conductivity2:standard_name = "sea_water_electrical_conductivity" ;
< 		conductivity2:units = "S m-1" ;
< 		conductivity2:coverage_content_type = "physicalMeasurement" ;
< 	double beam_transmission(depth) ;
< 		beam_transmission:_FillValue = NaN ;
< 		beam_transmission:long_name = "Percent of beam transmission of CTD measurement" ;
< 		beam_transmission:valid_max = 100. ;
< 		beam_transmission:valid_min = 0. ;
< 		beam_transmission:add_offset = 0. ;
< 		beam_transmission:scale_factor = 1. ;
< 		beam_transmission:standard_name = "volume_beam_attenuation_coefficient_of_radiative_flux_in_sea_water" ;
< 		beam_transmission:units = "%" ;
< 		beam_transmission:coverage_content_type = "physicalMeasurement" ;
< 	double fluorescence(depth) ;
< 		fluorescence:_FillValue = NaN ;
< 		fluorescence:long_name = "Fluorescence of CTD measurement" ;
< 		fluorescence:valid_max = 1.2009 ;
< 		fluorescence:valid_min = 0.8248 ;
< 		fluorescence:add_offset = 0. ;
< 		fluorescence:coordinates = "time depth latitude longitude" ;
< 		fluorescence:scale_factor = 1. ;
< 		fluorescence:standard_name = "fluorescence" ;
< 		fluorescence:units = "mg m-3" ;
< 		fluorescence:coverage_content_type = "physicalMeasurement" ;
< 	double par(depth) ;
< 		par:_FillValue = NaN ;
< 		par:long_name = "PAR of CTD measurement" ;
< 		par:valid_max = 1.e-12 ;
< 		par:valid_min = 1.e-12 ;
< 		par:add_offset = 0. ;
< 		par:coordinates = "time depth latitude longitude" ;
< 		par:scale_factor = 1. ;
< 		par:standard_name = "par" ;
< 		par:coverage_content_type = "physicalMeasurement" ;
< 	double salinity(depth) ;
< 		salinity:_FillValue = NaN ;
< 		salinity:long_name = "Salinity of CTD measurement" ;
< 		salinity:valid_max = 42. ;
< 		salinity:valid_min = 2. ;
< 		salinity:add_offset = 0. ;
< 		salinity:coordinates = "time depth latitude longitude" ;
< 		salinity:scale_factor = 1. ;
< 		salinity:standard_name = "sea_water_practical_salinity" ;
< 		salinity:units = "1" ;
< 		salinity:coverage_content_type = "physicalMeasurement" ;
< 	double salinity2(depth) ;
< 		salinity2:_FillValue = NaN ;
< 		salinity2:long_name = "Salinity of second CTD measurement" ;
< 		salinity2:valid_max = 42. ;
< 		salinity2:valid_min = 2. ;
< 		salinity2:add_offset = 0. ;
< 		salinity2:coordinates = "time depth latitude longitude" ;
< 		salinity2:scale_factor = 1. ;
< 		salinity2:standard_name = "sea_water_practical_salinity" ;
< 		salinity2:units = "1" ;
< 		salinity2:coverage_content_type = "physicalMeasurement" ;
< 	double potential_temperature(depth) ;
< 		potential_temperature:_FillValue = NaN ;
< 		potential_temperature:long_name = "Potential termperature of CTD measurement" ;
< 		potential_temperature:valid_max = 32. ;
< 		potential_temperature:valid_min = -1. ;
< 		potential_temperature:add_offset = 0. ;
< 		potential_temperature:coordinates = "time depth latitude longitude" ;
< 		potential_temperature:scale_factor = 1. ;
< 		potential_temperature:standard_name = "sea_water_potential_temperature" ;
< 		potential_temperature:units = "degrees_C" ;
< 		potential_temperature:coverage_content_type = "physicalMeasurement" ;
< 	double potential_temperature2(depth) ;
< 		potential_temperature2:_FillValue = NaN ;
< 		potential_temperature2:long_name = "Potential termperature of second CTD measurement" ;
< 		potential_temperature2:valid_max = 32. ;
< 		potential_temperature2:valid_min = -1. ;
< 		potential_temperature2:add_offset = 0. ;
< 		potential_temperature2:coordinates = "time depth latitude longitude" ;
< 		potential_temperature2:scale_factor = 1. ;
< 		potential_temperature2:standard_name = "sea_water_potential_temperature" ;
< 		potential_temperature2:units = "degrees_C" ;
< 		potential_temperature2:coverage_content_type = "physicalMeasurement" ;
< 	double density(depth) ;
< 		density:_FillValue = NaN ;
< 		density:long_name = "Density of CTD measurement" ;
< 		density:valid_max = 30. ;
< 		density:valid_min = 20. ;
< 		density:add_offset = 0. ;
< 		density:coordinates = "time depth latitude longitude" ;
< 		density:scale_factor = 1. ;
< 		density:standard_name = "sea_water_sigma_theta" ;
< 		density:units = "kg m-3" ;
< 		density:coverage_content_type = "physicalMeasurement" ;
< 	double density2(depth) ;
< 		density2:_FillValue = NaN ;
< 		density2:long_name = "Density of second CTD measurement" ;
< 		density2:valid_max = 30. ;
< 		density2:valid_min = 20. ;
< 		density2:add_offset = 0. ;
< 		density2:coordinates = "time depth latitude longitude" ;
< 		density2:scale_factor = 1. ;
< 		density2:standard_name = "sea_water_sigma_theta" ;
< 		density2:units = "kg m-3" ;
< 		density2:coverage_content_type = "physicalMeasurement" ;
< 	double oxygen(depth) ;
< 		oxygen:_FillValue = NaN ;
< 		oxygen:long_name = "Oxygen of CTD measurement" ;
< 		oxygen:valid_max = 7. ;
< 		oxygen:valid_min = 0. ;
< 		oxygen:add_offset = 0. ;
< 		oxygen:coordinates = "time depth latitude longitude" ;
< 		oxygen:scale_factor = 1. ;
< 		oxygen:standard_name = "volume_fraction_of_oxygen_in_sea_water" ;
< 		oxygen:units = "ml l-1" ;
< 		oxygen:coverage_content_type = "physicalMeasurement" ;
< 	double sound_velocity(depth) ;
< 		sound_velocity:_FillValue = NaN ;
< 		sound_velocity:long_name = "Sound velocity of CTD measurement" ;
< 		sound_velocity:valid_max = 1600. ;
< 		sound_velocity:valid_min = 1400. ;
< 		sound_velocity:add_offset = 0. ;
< 		sound_velocity:coordinates = "time depth latitude longitude" ;
< 		sound_velocity:scale_factor = 1. ;
< 		sound_velocity:standard_name = "speed_of_sound_in_sea_water" ;
< 		sound_velocity:units = "m s-1" ;
< 		sound_velocity:coverage_content_type = "physicalMeasurement" ;
< 	double sound_velocity2(depth) ;
< 		sound_velocity2:_FillValue = NaN ;
< 		sound_velocity2:long_name = "Sound velocity of second CTD measurement" ;
< 		sound_velocity2:valid_max = 1600. ;
< 		sound_velocity2:valid_min = 1400. ;
< 		sound_velocity2:add_offset = 0. ;
< 		sound_velocity2:coordinates = "time depth latitude longitude" ;
< 		sound_velocity2:scale_factor = 1. ;
< 		sound_velocity2:standard_name = "speed_of_sound_in_sea_water" ;
< 		sound_velocity2:units = "m s-1" ;
< 		sound_velocity2:coverage_content_type = "physicalMeasurement" ;
---
> 		depth:coverage_content_type = "referenceInformation" ;
> 
>     group: UnderwayCTD {
>         variables:
> 			double temperature(time) ;
> 				temperature:_FillValue = -9999. ;
> 				temperature:long_name = "Temperature of CTD measurement" ;
> 				temperature:valid_max = 32. ;
> 				temperature:valid_min = -1. ;
> 				temperature:coordinates = "time latitude longitude depth platform_id" ;
> 				temperature:standard_name = "sea_water_temperature" ;
> 				temperature:units = "degrees_C" ;
> 				temperature:coverage_content_type = "physicalMeasurement" ;
> 			double conductivity(time) ;
> 				conductivity:_FillValue = -9999. ;
> 				conductivity:long_name = "Conductivity of CTD measurement" ;
> 				conductivity:valid_max = 60. ;
> 				conductivity:valid_min = 0. ;
> 				conductivity:coordinates = "time latitude longitude depth platform_id" ;
> 				conductivity:standard_name = "sea_water_electrical_conductivity" ;
> 				conductivity:units = "S m-1" ;
> 				conductivity:coverage_content_type = "physicalMeasurement" ;
> 			double salinity(time) ;
> 				salinity:_FillValue = -9999. ;
> 				salinity:long_name = "Salinity of CTD measurement" ;
> 				salinity:valid_max = 42. ;
> 				salinity:valid_min = 2. ;
> 				salinity:coordinates = "time latitude longitude depth platform_id" ;
> 				salinity:standard_name = "sea_water_practical_salinity" ;
> 				salinity:units = "1" ;
> 				salinity:comments = "Salinity is assumed to be a ratio because of units=1. Provide more details about physical units in this field, e.g. (cm3 cm-3) for volumetric ratio." ;
> 				salinity:coverage_content_type = "physicalMeasurement" ;
> 			double density(time) ;
> 				density:_FillValue = -9999. ;
> 				density:long_name = "Density of CTD measurement" ;
> 				density:valid_max = 30. ;
> 				density:valid_min = 20. ;
> 				density:coordinates = "time latitude longitude depth platform_id" ;
> 				density:standard_name = "sea_water_sigma_theta" ;
> 				density:units = "kg m-3" ;
> 				density:coverage_content_type = "physicalMeasurement" ;
> 			double potential_temperature(time) ;
> 				potential_temperature:_FillValue = -9999. ;
> 				potential_temperature:long_name = "Potential termperature of CTD measurement" ;
> 				potential_temperature:valid_max = 32. ;
> 				potential_temperature:valid_min = -1. ;
> 				potential_temperature:coordinates = "time latitude longitude depth platform_id" ;
> 				potential_temperature:standard_name = "sea_water_potential_temperature" ;
> 				potential_temperature:units = "degrees_C" ;
> 				potential_temperature:coverage_content_type = "physicalMeasurement" ;
> 			double sound_velocity(time) ;
> 				sound_velocity:_FillValue = -9999. ;
> 				sound_velocity:long_name = "Sound velocity of CTD measurement" ;
> 				sound_velocity:valid_max = 1600. ;
> 				sound_velocity:valid_min = 1400. ;
> 				sound_velocity:coordinates = "time latitude longitude depth platform_id" ;
> 				sound_velocity:standard_name = "speed_of_sound_in_sea_water" ;
> 				sound_velocity:units = "m s-1" ;
> 				sound_velocity:coverage_content_type = "physicalMeasurement" ;
> 
> 		// group attributes:
> 		:description = "UnderwayCTD" ;
> 		:investigator = "Last Name, First Name" ;
> 		:instrument = "NULL" ;
> 		:platform = "NULL" ;
> 	}
> 
>     group: EcoCTD {
>         variables:
> 			double pressure(time) ;
> 				pressure:_FillValue = -9999. ;
> 				pressure:long_name = "Pressure of CTD measurement" ;
> 				pressure:valid_max = 1500. ;
> 				pressure:valid_min = -1. ;
> 				pressure:coordinates = "time depth latitude longitude platform_id" ;
> 				pressure:standard_name = "sea_water_pressure" ;
> 				pressure:units = "dbar" ;
> 				pressure:coverage_content_type = "physicalMeasurement" ;
> 			double temperature(time) ;
> 				temperature:_FillValue = -9999. ;
> 				temperature:long_name = "Temperature of second CTD measurement" ;
> 				temperature:valid_max = 32. ;
> 				temperature:valid_min = -1. ;
> 				temperature:coordinates = "time latitude longitude depth platform_id" ;
> 				temperature:standard_name = "sea_water_temperature" ;
> 				temperature:units = "degrees_C" ;
> 				temperature:coverage_content_type = "physicalMeasurement" ;
> 			double conductivity(time) ;
> 				conductivity:_FillValue = -9999. ;
> 				conductivity:long_name = "Conductivity of second CTD measurement" ;
> 				conductivity:valid_max = 60. ;
> 				conductivity:valid_min = 0. ;
> 				conductivity:coordinates = "time latitude longitude depth platform_id" ;
> 				conductivity:standard_name = "sea_water_electrical_conductivity" ;
> 				conductivity:units = "S m-1" ;
> 				conductivity:coverage_content_type = "physicalMeasurement" ;
> 			double salinity(time) ;
> 				salinity:_FillValue = -9999. ;
> 				salinity:long_name = "Salinity of second CTD measurement" ;
> 				salinity:valid_max = 42. ;
> 				salinity:valid_min = 2. ;
> 				salinity:coordinates = "time latitude longitude depth platform_id" ;
> 				salinity:standard_name = "sea_water_practical_salinity" ;
> 				salinity:units = "1" ;
> 				salinity:comments = "Salinity is assumed to be a ratio because of units=1. Provide more details about physical units in this field, e.g. (cm3 cm-3) for volumetric ratio." ;
> 				salinity:coverage_content_type = "physicalMeasurement" ;
> 			double potential_temperature(time) ;
> 				potential_temperature:_FillValue = -9999. ;
> 				potential_temperature:long_name = "Potential termperature of second CTD measurement" ;
> 				potential_temperature:valid_max = 32. ;
> 				potential_temperature:valid_min = -1. ;
> 				potential_temperature:coordinates = "time latitude longitude depth platform_id" ;
> 				potential_temperature:standard_name = "sea_water_potential_temperature" ;
> 				potential_temperature:units = "degrees_C" ;
> 				potential_temperature:coverage_content_type = "physicalMeasurement" ;
> 			double sound_velocity(time) ;
> 				sound_velocity:_FillValue = -9999. ;
> 				sound_velocity:long_name = "Sound velocity of second CTD measurement" ;
> 				sound_velocity:valid_max = 1600. ;
> 				sound_velocity:valid_min = 1400. ;
> 				sound_velocity:coordinates = "time latitude longitude depth platform_id" ;
> 				sound_velocity:standard_name = "speed_of_sound_in_sea_water" ;
> 				sound_velocity:units = "m s-1" ;
> 				sound_velocity:coverage_content_type = "physicalMeasurement" ;
> 			double density(time) ;
> 				density:_FillValue = -9999. ;
> 				density:long_name = "Density of second CTD measurement" ;
> 				density:valid_max = 30. ;
> 				density:valid_min = 20. ;
> 				density:coordinates = "time latitude longitude depth platform_id" ;
> 				density:standard_name = "sea_water_sigma_theta" ;
> 				density:units = "kg m-3" ;
> 				density:coverage_content_type = "physicalMeasurement" ;
> 			double beam_transmission(time) ;
> 				beam_transmission:_FillValue = -9999. ;
> 				beam_transmission:long_name = "Percent of beam transmission of CTD measurement" ;
> 				beam_transmission:valid_max = 100. ;
> 				beam_transmission:valid_min = 0. ;
> 				beam_transmission:standard_name = "volume_beam_attenuation_coefficient_of_radiative_flux_in_sea_water" ;
> 				beam_transmission:units = "%" ;
> 				beam_transmission:coverage_content_type = "physicalMeasurement" ;
> 			double fluorescence(time) ;
> 				fluorescence:_FillValue = -9999. ;
> 				fluorescence:long_name = "Fluorescence of CTD measurement" ;
> 				fluorescence:valid_max = 1.2009 ;
> 				fluorescence:valid_min = 0.8248 ;
> 				fluorescence:coordinates = "time latitude longitude depth platform_id" ;
> 				fluorescence:standard_name = "fluorescence" ;
> 				fluorescence:units = "mg m-3" ;
> 				fluorescence:coverage_content_type = "physicalMeasurement" ;
> 			double par(time) ;
> 				par:_FillValue = -9999. ;
> 				par:long_name = "PAR of CTD measurement" ;
> 				par:valid_max = 1.e-12 ;
> 				par:valid_min = 1.e-12 ;
> 				par:coordinates = "time latitude longitude depth platform_id" ;
> 				par:standard_name = "par" ;
> 				par:coverage_content_type = "physicalMeasurement" ;
> 			double oxygen(time) ;
> 				oxygen:_FillValue = -9999. ;
> 				oxygen:long_name = "Oxygen of CTD measurement" ;
> 				oxygen:valid_max = 7. ;
> 				oxygen:valid_min = 0. ;
> 				oxygen:coordinates = "time latitude longitude depth platform_id" ;
> 				oxygen:standard_name = "volume_fraction_of_oxygen_in_sea_water" ;
> 				oxygen:units = "ml l-1" ;
> 				oxygen:coverage_content_type = "physicalMeasurement" ;
> 
> 		// group attributes:
> 		:description = "EcoCTD";
> 		:investigator = "Last Name, First Name" ;
> 		:instrument = "NULL" ;
> 		:platform = "NULL" ;
> 	}
