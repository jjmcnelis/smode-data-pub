netcdf S-MODE_PFC_seaglider_\#\# {
dimensions:
	ctd_time = 864583 ;
	dive = 820 ;
variables:
	double ctd_depth(ctd_time) ;
		ctd_depth:_FillValue = NaN ;
		ctd_depth:long_name = "Depth" ;
		ctd_depth:valid_max = 2000. ;
		ctd_depth:valid_min = 0. ;
		ctd_depth:axis = "Z" ;
		ctd_depth:positive = "down" ;
		ctd_depth:standard_name = "depth" ;
		ctd_depth:units = "m" ;
		ctd_depth:coverage_content_type = "coordinate" ;
	double ctd_data_point_dive_number(ctd_time) ;
		ctd_data_point_dive_number:_FillValue = -2147483648. ;
		ctd_data_point_dive_number:long_name = "Dive Number for given ctd_data_point observation" ;
		ctd_data_point_dive_number:add_offset = 0. ;
		ctd_data_point_dive_number:scale_factor = 1. ;
		ctd_data_point_dive_number:comment = "Dive number for given ctd_data_point observation" ;
		ctd_data_point_dive_number:coordinates = "ctd_time longitude latitude ctd_depth" ;
	double ctd_time(ctd_time) ;
		ctd_time:long_name = "Time of CTD sample" ;
		ctd_time:axis = "T" ;
		ctd_time:standard_name = "time" ;
		ctd_time:units = "days since 1950-01-01T00:00:00" ;
		ctd_time:coverage_content_type = "coordinate" ;
	double longitude(ctd_time) ;
		longitude:_FillValue = NaN ;
		longitude:long_name = "Longitude of the sample based on hdm DAC" ;
		longitude:valid_max = 180. ;
		longitude:valid_min = -180. ;
		longitude:axis = "X" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "coordinate" ;
	double latitude(ctd_time) ;
		latitude:_FillValue = NaN ;
		latitude:long_name = "Latitude of the sample based on hdm DAC" ;
		latitude:valid_max = 90. ;
		latitude:valid_min = -90. ;
		latitude:axis = "Y" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "coordinate" ;
	double conductivity(ctd_time) ;
		conductivity:_FillValue = NaN ;
		conductivity:long_name = "Conductivity corrected for anomalies" ;
		conductivity:valid_max = 60. ;
		conductivity:valid_min = 0. ;
		conductivity:add_offset = 0. ;
		conductivity:scale_factor = 1. ;
		conductivity:standard_name = "sea_water_electrical_conductivity" ;
		conductivity:units = "S m-1" ;
		conductivity:coordinates = "ctd_time longitude latitude ctd_depth" ;
		conductivity:coverage_content_type = "physicalMeasurement" ;
	double ctd_pressure(ctd_time) ;
		ctd_pressure:_FillValue = NaN ;
		ctd_pressure:long_name = "Pressure at CTD thermistor" ;
		ctd_pressure:valid_max = 2000. ;
		ctd_pressure:valid_min = -1. ;
		ctd_pressure:add_offset = 0. ;
		ctd_pressure:scale_factor = 1. ;
		ctd_pressure:standard_name = "sea_water_pressure" ;
		ctd_pressure:units = "dbar" ;
		ctd_pressure:coordinates = "ctd_time longitude latitude ctd_depth" ;
		ctd_pressure:coverage_content_type = "physicalMeasurement" ;
	double temperature(ctd_time) ;
		temperature:_FillValue = NaN ;
		temperature:long_name = "Temperature (in situ) corrected for thermistor first-order lag" ;
		temperature:valid_max = 32. ;
		temperature:valid_min = -1. ;
		temperature:add_offset = 0. ;
		temperature:scale_factor = 1. ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "degrees_C" ;
		temperature:coordinates = "ctd_time longitude latitude ctd_depth" ;
		temperature:coverage_content_type = "physicalMeasurement" ;
	double salinity(ctd_time) ;
		salinity:_FillValue = NaN ;
		salinity:long_name = "Salinity corrected for thermal-inertia effects (PSU)" ;
		salinity:valid_max = 42. ;
		salinity:valid_min = 2. ;
		salinity:add_offset = 0. ;
		salinity:scale_factor = 1. ;
		salinity:standard_name = "sea_water_practical_salinity" ;
		salinity:units = "1" ;
		salinity:coordinates = "ctd_time longitude latitude ctd_depth" ;
		salinity:coverage_content_type = "physicalMeasurement" ;
	double mean_time(dive) ;
		mean_time:long_name = "Mean time of the dive" ;
		mean_time:standard_name = "time" ;
		mean_time:units = "days since 1950-01-01T00:00:00" ;
		mean_time:coverage_content_type = "coordinate" ;
	double mean_longitude(dive) ;
		mean_longitude:_FillValue = NaN ;
		mean_longitude:long_name = "Mean longitude of the dive" ;
		mean_longitude:valid_max = 180. ;
		mean_longitude:valid_min = -180. ;
		mean_longitude:standard_name = "longitude" ;
		mean_longitude:units = "degrees_east" ;
		mean_longitude:coverage_content_type = "coordinate" ;
	double mean_latitude(dive) ;
		mean_latitude:_FillValue = NaN ;
		mean_latitude:long_name = "Mean latitude of the dive" ;
		mean_latitude:valid_max = 90. ;
		mean_latitude:valid_min = -90. ;
		mean_latitude:standard_name = "latitude" ;
		mean_latitude:units = "degrees_north" ;
		mean_latitude:coverage_content_type = "coordinate" ;
	double start_time(dive) ;
		start_time:long_name = "Starting time of the dive" ;
		start_time:standard_name = "time" ;
		start_time:units = "days since 1950-01-01T00:00:00" ;
		start_time:coverage_content_type = "coordinate" ;
	double start_longitude(dive) ;
		start_longitude:_FillValue = NaN ;
		start_longitude:long_name = "Starting longitude of the dive" ;
		start_longitude:valid_max = 180. ;
		start_longitude:valid_min = -180. ;
		start_longitude:standard_name = "longitude" ;
		start_longitude:units = "degrees_east" ;
		start_longitude:coverage_content_type = "coordinate" ;
	double start_latitude(dive) ;
		start_latitude:_FillValue = NaN ;
		start_latitude:long_name = "Starting latitude of the dive" ;
		start_latitude:valid_max = 90. ;
		start_latitude:valid_min = -90. ;
		start_latitude:standard_name = "latitude" ;
		start_latitude:units = "degrees_north" ;
		start_latitude:coverage_content_type = "coordinate" ;
	double end_time(dive) ;
		end_time:long_name = "Ending time of the dive" ;
		end_time:standard_name = "time" ;
		end_time:units = "days since 1950-01-01T00:00:00" ;
		end_time:coverage_content_type = "coordinate" ;
	double end_longitude(dive) ;
		end_longitude:_FillValue = NaN ;
		end_longitude:long_name = "Ending longitude of the dive" ;
		end_longitude:valid_max = 180. ;
		end_longitude:valid_min = -180. ;
		end_longitude:standard_name = "longitude" ;
		end_longitude:units = "degrees_east" ;
		end_longitude:coverage_content_type = "coordinate" ;
	double end_latitude(dive) ;
		end_latitude:_FillValue = NaN ;
		end_latitude:long_name = "Ending latitude of the dive" ;
		end_latitude:valid_max = 90. ;
		end_latitude:valid_min = -90. ;
		end_latitude:standard_name = "latitude" ;
		end_latitude:units = "degrees_north" ;
		end_latitude:coverage_content_type = "coordinate" ;

// global attributes:
		:DOI = "10.5067/SMODE-GLID1" ;
		:title = "S-MODE  Pilot Field Campaign Fall 2020 Temperature and Salinity from Seagliders<, XXXX>" ;
		:summary = "S-MODE  Pilot Field Campaign Fall 2020 Temperature and Salinity from Seagliders<, XXXX>" ;
		:keywords = "EARTH SCIENCE > OCEANS > SALINITY/DENSITY > CONDUCTIVITY, EARTH SCIENCE > OCEANS > OCEAN TEMPERATURE > TEMPERATURE PROFILES, EARTH SCIENCE > OCEANS > SALINITY/DENSITY > SALINITY" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:conventions = "CF-1.8, ACDD-1.3" ;
		:id = "PO.DAAC-SMODE-GLID1" ;
		:uuid = "784c15f0-1a8e-49ad-9d48-653066dc2450" ;
		:naming_authority = "gov.nasa" ;
		:featureType = "trajectory" ;
		:cdm_data_type = "Trajectory" ;
		:source = "TBD" ;
		:platform = "In Situ Ocean-based Platforms > > SEAGLIDER" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:instrument = "In Situ/Laboratory Instruments > Profilers/Sounders > > > CTD" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:processing_level = "L2" ;
		:standard_name_vocabulary = "CF Standard Name Table v72" ;
		:acknowledgement = "TBD" ;
		:comment = "" ;
		:license = "S-MODE data are considered experimental and not to be used for any purpose for which life or property is potentially at risk. Distributor assumes no responsibility for the manner in which the data are used. Otherwise data are free for public use." ;
		:product_version = "1" ;
		:metadata_link = "https://doi.org/10.5067/SMODE-GLID1" ;
		:creator_name = "Tom Farrar" ;
		:creator_email = "jfarrar@whoi.edu" ;
		:creator_type = "person" ;
		:creator_institution = "WHOI/" ;
		:institution = "WHOI/" ;
		:project = "Sub-Mesoscale Ocean Dynamics Experiment (S-MODE)" ;
		:program = "NASA Earth Venture Suborbital-3 (EVS-3)" ;
		:contributor_name = "Frederick Bingham" ;
		:contributor_role = "Project Data Manager" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center, Jet Propulsion Laboratory, NASA" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:sea_name = "Pacific" ;
		:geospatial_lat_min = 8.99499833333333 ;
		:geospatial_lat_max = 12.0227483333333 ;
		:geospatial_lat_units = "degrees" ;
		:geospatial_lat_resolution = "0.1" ;
		:geospatial_lon_min = -126.62557 ;
		:geospatial_lon_max = -122.12858 ;
		:geospatial_lon_units = "degrees" ;
		:geospatial_lon_resolution = "0.1" ;
		:geospatial_vertical_min = 8.37780569335051e-05 ;
		:geospatial_vertical_max = 1001.54380074156 ;
		:geospatial_vertical_resolution = "1" ;
		:geospatial_vertical_units = "m" ;
		:geospatial_vertical_positive = "down" ;
		:time_coverage_start = "26-Aug-2016 15:49:21" ;
		:time_coverage_end = "08-May-2017 17:16:34" ;
		:date_created = "01-Sep-2020 14:14:02" ;
}
