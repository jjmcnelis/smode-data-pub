netcdf S-MODE_PFC_OC2004B_rawinsonde_\#\# {
dimensions:
	profile_time = 82 ;
	nz = 20000 ;
variables:
	double profile_time(profile_time) ;
		profile_time:long_name = "Profile Time of Rawinsonde" ;
		profile_time:axis = "T" ;
		profile_time:standard_name = "time" ;
		profile_time:units = "days since 1950-01-01T00:00:00" ;
		profile_time:coverage_content_type = "coordinate" ;
	double profile_longitude(profile_time) ;
		profile_longitude:_FillValue = NaN ;
		profile_longitude:long_name = "Profile Longitude of Rawinsonde" ;
		profile_longitude:valid_max = 180. ;
		profile_longitude:valid_min = -180. ;
		profile_longitude:standard_name = "longitude" ;
		profile_longitude:units = "degrees_east" ;
		profile_longitude:coverage_content_type = "coordinate" ;
	double profile_latitude(profile_time) ;
		profile_latitude:_FillValue = NaN ;
		profile_latitude:long_name = "Profile Latitude of Rawinsonde" ;
		profile_latitude:valid_max = 90. ;
		profile_latitude:valid_min = -90. ;
		profile_latitude:standard_name = "latitude" ;
		profile_latitude:units = "degrees_north" ;
		profile_latitude:coverage_content_type = "coordinate" ;
	double time(profile_time, nz) ;
		time:long_name = "Time of Rawinsonde" ;
		time:standard_name = "time" ;
		time:units = "days since 1950-01-01T00:00:00" ;
		time:coverage_content_type = "coordinate" ;
	double longitude(profile_time, nz) ;
		longitude:_FillValue = NaN ;
		longitude:long_name = "Longitude of Rawinsonde" ;
		longitude:valid_max = 180. ;
		longitude:valid_min = -180. ;
		longitude:axis = "X" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "coordinate" ;
	double latitude(profile_time, nz) ;
		latitude:_FillValue = NaN ;
		latitude:long_name = "Latitude of Rawinsonde" ;
		latitude:valid_max = 90. ;
		latitude:valid_min = -90. ;
		latitude:axis = "Y" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "coordinate" ;
	double altitude(profile_time, nz) ;
		altitude:_FillValue = NaN ;
		altitude:long_name = "GPS Altitude above MSL" ;
		altitude:valid_max = 20000. ;
		altitude:valid_min = 0. ;
		altitude:axis = "Z" ;
		altitude:positive = "up" ;
		altitude:standard_name = "altitude" ;
		altitude:units = "m" ;
		altitude:coverage_content_type = "coordinate" ;
	double air_pressure(profile_time, nz) ;
		air_pressure:_FillValue = NaN ;
		air_pressure:long_name = "Air Pressure" ;
		air_pressure:valid_max = 1021. ;
		air_pressure:valid_min = 12.3934488 ;
		air_pressure:add_offset = "0" ;
		air_pressure:scale_factor = 1. ;
		air_pressure:standard_name = "air_pressure" ;
		air_pressure:units = "mbar" ;
		air_pressure:coordinates = "profile_time altitude latitude longitude" ;
		air_pressure:coverage_content_type = "physicalMeasurement" ;
	double air_temperature(profile_time, nz) ;
		air_temperature:_FillValue = NaN ;
		air_temperature:long_name = "Air Temperature" ;
		air_temperature:valid_max = 29.0737999999999 ;
		air_temperature:valid_min = -85.9452 ;
		air_temperature:add_offset = "0" ;
		air_temperature:scale_factor = 1. ;
		air_temperature:standard_name = "air_temperature" ;
		air_temperature:units = "degrees_C" ;
		air_temperature:coordinates = "profile_time altitude latitude longitude" ;
		air_temperature:coverage_content_type = "physicalMeasurement" ;
	double relative_humidity(profile_time, nz) ;
		relative_humidity:_FillValue = NaN ;
		relative_humidity:long_name = "Relative Humidity" ;
		relative_humidity:valid_max = 100. ;
		relative_humidity:valid_min = 0. ;
		relative_humidity:add_offset = "0" ;
		relative_humidity:scale_factor = 1. ;
		relative_humidity:standard_name = "relative_humidity" ;
		relative_humidity:units = "%" ;
		relative_humidity:coordinates = "profile_time altitude latitude longitude" ;
		relative_humidity:coverage_content_type = "physicalMeasurement" ;
	double wind_direction(profile_time, nz) ;
		wind_direction:_FillValue = NaN ;
		wind_direction:long_name = "Wind Direction" ;
		wind_direction:valid_max = 360. ;
		wind_direction:valid_min = 0. ;
		wind_direction:add_offset = "0" ;
		wind_direction:scale_factor = 1. ;
		wind_direction:standard_name = "wind_from_direction" ;
		wind_direction:units = "degrees" ;
		wind_direction:coordinates = "profile_time altitude latitude longitude" ;
		wind_direction:coverage_content_type = "physicalMeasurement" ;
	double wind_speed(profile_time, nz) ;
		wind_speed:_FillValue = NaN ;
		wind_speed:long_name = "Wind Speed" ;
		wind_speed:valid_max = 40. ;
		wind_speed:valid_min = 0. ;
		wind_speed:add_offset = "0" ;
		wind_speed:scale_factor = 1. ;
		wind_speed:standard_name = "wind_speed" ;
		wind_speed:units = "m s-1" ;
		wind_speed:coordinates = "profile_time altitude latitude longitude" ;
		wind_speed:coverage_content_type = "physicalMeasurement" ;
	double eastward_wind_component(profile_time, nz) ;
		eastward_wind_component:_FillValue = NaN ;
		eastward_wind_component:long_name = "Eastward Wind Component" ;
		eastward_wind_component:valid_max = 40. ;
		eastward_wind_component:valid_min = -40. ;
		eastward_wind_component:add_offset = "0" ;
		eastward_wind_component:scale_factor = 1. ;
		eastward_wind_component:standard_name = "eastward_wind" ;
		eastward_wind_component:units = "m s-1" ;
		eastward_wind_component:coordinates = "profile_time altitude latitude longitude" ;
		eastward_wind_component:coverage_content_type = "physicalMeasurement" ;
	double northward_wind_component(profile_time, nz) ;
		northward_wind_component:_FillValue = NaN ;
		northward_wind_component:long_name = "Northward Wind Component" ;
		northward_wind_component:valid_max = 40. ;
		northward_wind_component:valid_min = -40. ;
		northward_wind_component:add_offset = "0" ;
		northward_wind_component:scale_factor = 1. ;
		northward_wind_component:standard_name = "northward_wind" ;
		northward_wind_component:units = "m s-1" ;
		northward_wind_component:coordinates = "profile_time altitude latitude longitude" ;
		northward_wind_component:coverage_content_type = "physicalMeasurement" ;

// global attributes:
		:DOI = "10.5067/SMODE-SONDE" ;
		:title = "S-MODE  Pilot Field Campaign Fall 2020 Meteorological Data from Rawinsondes deployed by R/V Oceanus<, XXXX>" ;
		:summary = "S-MODE  Pilot Field Campaign Fall 2020 Meteorological Data from Rawinsondes deployed by R/V Oceanus<, XXXX>" ;
		:keywords = "EARTH SCIENCE > ATMOSPHERE > ATMOSPHERIC WINDS > WIND PROFILES, EARTH SCIENCE > OCEANS > OCEAN WINDS > SURFACE WINDS, EARTH SCIENCE > ATMOSPHERE > ATMOSPHERIC TEMPERATURE > AIR TEMPERATURE, EARTH SCIENCE > ATMOSPHERE > HUMIDITY INDICES > HUMIDITY, EARTH SCIENCE > ATMOSPHERE > ATMOSPHERIC PRESSURE > ATMOSPHERIC PRESSURE MEASUREMENTS" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:conventions = "CF-1.8, ACDD-1.3" ;
		:id = "PO.DAAC-SMODE-SONDE" ;
		:uuid = "4e368f4e-1648-4260-8bc0-5903523cb27e" ;
		:naming_authority = "gov.nasa" ;
		:featureType = "profile" ;
		:cdm_data_type = "Station" ;
		:source = "TBD" ;
		:platform = "In Situ Ocean-based Platforms > SHIPS > RV Oceanus, Balloons/Rockets > > RAWINSONDES, Balloons/Rockets > > RADIOSONDES" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:instrument = "Earth Remote Sensing Instruments > Passive Remote Sensing > Profilers/Sounders > > RADIOSONDES" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:processing_level = "L2" ;
		:standard_name_vocabulary = "CF Standard Name Table v72" ;
		:acknowledgement = "TBD" ;
		:comment = "" ;
		:license = "S-MODE data are considered experimental and not to be used for any purpose for which life or property is potentially at risk. Distributor assumes no responsibility for the manner in which the data are used. Otherwise data are free for public use." ;
		:product_version = "1" ;
		:metadata_link = "https://doi.org/10.5067/SMODE-SONDE" ;
		:creator_name = "Larry O\'Neill" ;
		:creator_email = "loneill@coas.oregonstate.edu" ;
		:creator_type = "person" ;
		:creator_institution = "OR-STATE/" ;
		:institution = "OR-STATE/" ;
		:project = "Sub-Mesoscale Ocean Dynamics Experiment (S-MODE)" ;
		:program = "NASA Earth Venture Suborbital-3 (EVS-3)" ;
		:contributor_name = "Frederick Bingham" ;
		:contributor_role = "Project Data Manager" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center, Jet Propulsion Laboratory, NASA" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:sea_name = "Pacific" ;
		:geospatial_lat_min = 5.03647267240922 ;
		:geospatial_lat_max = 13.5394171775961 ;
		:geospatial_lat_units = "degrees" ;
		:geospatial_lat_resolution = "0.1" ;
		:geospatial_lon_min = -133.216191968924 ;
		:geospatial_lon_max = -123.322785250482 ;
		:geospatial_lon_units = "degrees" ;
		:geospatial_lon_resolution = "0.1" ;
		:geospatial_vertical_min = 2.99196165357995 ;
		:geospatial_vertical_max = 29544.1579589844 ;
		:geospatial_vertical_resolution = "1" ;
		:geospatial_vertical_units = "m" ;
		:geospatial_vertical_positive = "up" ;
		:time_coverage_start = "20-Aug-2016 01:56:45" ;
		:time_coverage_end = "14-Sep-2016 17:36:26" ;
		:date_created = "01-Sep-2020 14:12:34" ;
}
