netcdf S-MODE_PFC_OC2004B_ctd_\#\# {
dimensions:
	time = 1 ;
	depth = 79246 ;
variables:
	double time(time) ;
		time:long_name = "Time of CTD measurement" ;
		time:axis = "T" ;
		time:standard_name = "time" ;
		time:units = "days since 1950-01-01T00:00:00" ;
		time:coverage_content_type = "coordinate" ;
	double latitude(time) ;
		latitude:_FillValue = NaN ;
		latitude:long_name = "Latitude of CTD measurement" ;
		latitude:valid_max = 90. ;
		latitude:valid_min = -90. ;
		latitude:axis = "Y" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "coordinate" ;
	double longitude(time) ;
		longitude:_FillValue = NaN ;
		longitude:long_name = "Longitude of CTD measurement" ;
		longitude:valid_max = 180. ;
		longitude:valid_min = -180. ;
		longitude:axis = "X" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "coordinate" ;
	double depth(depth) ;
		depth:_FillValue = NaN ;
		depth:long_name = "Depth of CTD measurement" ;
		depth:valid_max = 1500. ;
		depth:valid_min = 0. ;
		depth:axis = "Z" ;
		depth:positive = "down" ;
		depth:standard_name = "depth" ;
		depth:units = "m" ;
		depth:coverage_content_type = "coordinate" ;
	double pressure(depth) ;
		pressure:_FillValue = NaN ;
		pressure:long_name = "Pressure of CTD measurement" ;
		pressure:valid_max = 1500. ;
		pressure:valid_min = -1. ;
		pressure:add_offset = 0. ;
		pressure:coordinates = "time depth latitude longitude" ;
		pressure:scale_factor = 1. ;
		pressure:standard_name = "sea_water_pressure" ;
		pressure:units = "dbar" ;
		pressure:coverage_content_type = "physicalMeasurement" ;
	double temperature(depth) ;
		temperature:_FillValue = NaN ;
		temperature:long_name = "Temperature of CTD measurement" ;
		temperature:valid_max = 32. ;
		temperature:valid_min = -1. ;
		temperature:add_offset = 0. ;
		temperature:coordinates = "time depth latitude longitude" ;
		temperature:scale_factor = 1. ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "degrees_C" ;
		temperature:coverage_content_type = "physicalMeasurement" ;
	double temperature2(depth) ;
		temperature2:_FillValue = NaN ;
		temperature2:long_name = "Temperature of second CTD measurement" ;
		temperature2:valid_max = 32. ;
		temperature2:valid_min = -1. ;
		temperature2:add_offset = 0. ;
		temperature2:coordinates = "time depth latitude longitude" ;
		temperature2:scale_factor = 1. ;
		temperature2:standard_name = "sea_water_temperature" ;
		temperature2:units = "degrees_C" ;
		temperature2:coverage_content_type = "physicalMeasurement" ;
	double conductivity(depth) ;
		conductivity:_FillValue = NaN ;
		conductivity:long_name = "Conductivity of CTD measurement" ;
		conductivity:valid_max = 60. ;
		conductivity:valid_min = 0. ;
		conductivity:add_offset = 0. ;
		conductivity:coordinates = "time depth latitude longitude" ;
		conductivity:scale_factor = 1. ;
		conductivity:standard_name = "sea_water_electrical_conductivity" ;
		conductivity:units = "S m-1" ;
		conductivity:coverage_content_type = "physicalMeasurement" ;
	double conductivity2(depth) ;
		conductivity2:_FillValue = NaN ;
		conductivity2:long_name = "Conductivity of second CTD measurement" ;
		conductivity2:valid_max = 60. ;
		conductivity2:valid_min = 0. ;
		conductivity2:add_offset = 0. ;
		conductivity2:coordinates = "time depth latitude longitude" ;
		conductivity2:scale_factor = 1. ;
		conductivity2:standard_name = "sea_water_electrical_conductivity" ;
		conductivity2:units = "S m-1" ;
		conductivity2:coverage_content_type = "physicalMeasurement" ;
	double beam_transmission(depth) ;
		beam_transmission:_FillValue = NaN ;
		beam_transmission:long_name = "Percent of beam transmission of CTD measurement" ;
		beam_transmission:valid_max = 100. ;
		beam_transmission:valid_min = 0. ;
		beam_transmission:add_offset = 0. ;
		beam_transmission:scale_factor = 1. ;
		beam_transmission:standard_name = "volume_beam_attenuation_coefficient_of_radiative_flux_in_sea_water" ;
		beam_transmission:units = "%" ;
		beam_transmission:coverage_content_type = "physicalMeasurement" ;
	double fluorescence(depth) ;
		fluorescence:_FillValue = NaN ;
		fluorescence:long_name = "Fluorescence of CTD measurement" ;
		fluorescence:valid_max = 1.2009 ;
		fluorescence:valid_min = 0.8248 ;
		fluorescence:add_offset = 0. ;
		fluorescence:coordinates = "time depth latitude longitude" ;
		fluorescence:scale_factor = 1. ;
		fluorescence:standard_name = "fluorescence" ;
		fluorescence:units = "mg m-3" ;
		fluorescence:coverage_content_type = "physicalMeasurement" ;
	double par(depth) ;
		par:_FillValue = NaN ;
		par:long_name = "PAR of CTD measurement" ;
		par:valid_max = 1.e-12 ;
		par:valid_min = 1.e-12 ;
		par:add_offset = 0. ;
		par:coordinates = "time depth latitude longitude" ;
		par:scale_factor = 1. ;
		par:standard_name = "par" ;
		par:coverage_content_type = "physicalMeasurement" ;
	double salinity(depth) ;
		salinity:_FillValue = NaN ;
		salinity:long_name = "Salinity of CTD measurement" ;
		salinity:valid_max = 42. ;
		salinity:valid_min = 2. ;
		salinity:add_offset = 0. ;
		salinity:coordinates = "time depth latitude longitude" ;
		salinity:scale_factor = 1. ;
		salinity:standard_name = "sea_water_practical_salinity" ;
		salinity:units = "1" ;
		salinity:coverage_content_type = "physicalMeasurement" ;
	double salinity2(depth) ;
		salinity2:_FillValue = NaN ;
		salinity2:long_name = "Salinity of second CTD measurement" ;
		salinity2:valid_max = 42. ;
		salinity2:valid_min = 2. ;
		salinity2:add_offset = 0. ;
		salinity2:coordinates = "time depth latitude longitude" ;
		salinity2:scale_factor = 1. ;
		salinity2:standard_name = "sea_water_practical_salinity" ;
		salinity2:units = "1" ;
		salinity2:coverage_content_type = "physicalMeasurement" ;
	double potential_temperature(depth) ;
		potential_temperature:_FillValue = NaN ;
		potential_temperature:long_name = "Potential termperature of CTD measurement" ;
		potential_temperature:valid_max = 32. ;
		potential_temperature:valid_min = -1. ;
		potential_temperature:add_offset = 0. ;
		potential_temperature:coordinates = "time depth latitude longitude" ;
		potential_temperature:scale_factor = 1. ;
		potential_temperature:standard_name = "sea_water_potential_temperature" ;
		potential_temperature:units = "degrees_C" ;
		potential_temperature:coverage_content_type = "physicalMeasurement" ;
	double potential_temperature2(depth) ;
		potential_temperature2:_FillValue = NaN ;
		potential_temperature2:long_name = "Potential termperature of second CTD measurement" ;
		potential_temperature2:valid_max = 32. ;
		potential_temperature2:valid_min = -1. ;
		potential_temperature2:add_offset = 0. ;
		potential_temperature2:coordinates = "time depth latitude longitude" ;
		potential_temperature2:scale_factor = 1. ;
		potential_temperature2:standard_name = "sea_water_potential_temperature" ;
		potential_temperature2:units = "degrees_C" ;
		potential_temperature2:coverage_content_type = "physicalMeasurement" ;
	double density(depth) ;
		density:_FillValue = NaN ;
		density:long_name = "Density of CTD measurement" ;
		density:valid_max = 30. ;
		density:valid_min = 20. ;
		density:add_offset = 0. ;
		density:coordinates = "time depth latitude longitude" ;
		density:scale_factor = 1. ;
		density:standard_name = "sea_water_sigma_theta" ;
		density:units = "kg m-3" ;
		density:coverage_content_type = "physicalMeasurement" ;
	double density2(depth) ;
		density2:_FillValue = NaN ;
		density2:long_name = "Density of second CTD measurement" ;
		density2:valid_max = 30. ;
		density2:valid_min = 20. ;
		density2:add_offset = 0. ;
		density2:coordinates = "time depth latitude longitude" ;
		density2:scale_factor = 1. ;
		density2:standard_name = "sea_water_sigma_theta" ;
		density2:units = "kg m-3" ;
		density2:coverage_content_type = "physicalMeasurement" ;
	double oxygen(depth) ;
		oxygen:_FillValue = NaN ;
		oxygen:long_name = "Oxygen of CTD measurement" ;
		oxygen:valid_max = 7. ;
		oxygen:valid_min = 0. ;
		oxygen:add_offset = 0. ;
		oxygen:coordinates = "time depth latitude longitude" ;
		oxygen:scale_factor = 1. ;
		oxygen:standard_name = "volume_fraction_of_oxygen_in_sea_water" ;
		oxygen:units = "ml l-1" ;
		oxygen:coverage_content_type = "physicalMeasurement" ;
	double sound_velocity(depth) ;
		sound_velocity:_FillValue = NaN ;
		sound_velocity:long_name = "Sound velocity of CTD measurement" ;
		sound_velocity:valid_max = 1600. ;
		sound_velocity:valid_min = 1400. ;
		sound_velocity:add_offset = 0. ;
		sound_velocity:coordinates = "time depth latitude longitude" ;
		sound_velocity:scale_factor = 1. ;
		sound_velocity:standard_name = "speed_of_sound_in_sea_water" ;
		sound_velocity:units = "m s-1" ;
		sound_velocity:coverage_content_type = "physicalMeasurement" ;
	double sound_velocity2(depth) ;
		sound_velocity2:_FillValue = NaN ;
		sound_velocity2:long_name = "Sound velocity of second CTD measurement" ;
		sound_velocity2:valid_max = 1600. ;
		sound_velocity2:valid_min = 1400. ;
		sound_velocity2:add_offset = 0. ;
		sound_velocity2:coordinates = "time depth latitude longitude" ;
		sound_velocity2:scale_factor = 1. ;
		sound_velocity2:standard_name = "speed_of_sound_in_sea_water" ;
		sound_velocity2:units = "m s-1" ;
		sound_velocity2:coverage_content_type = "physicalMeasurement" ;

// global attributes:
		:DOI = "10.5067/SMODE-RVCTD" ;
		:title = "S-MODE Pilot Field Campaign Fall 2020 Shipboard CTD measurements from the R/V Oceanus<, XXXX>" ;
		:summary = "S-MODE Pilot Field Campaign Fall 2020 Shipboard CTD measurements from the R/V Oceanus<, XXXX>" ;
		:keywords = "EARTH SCIENCE > OCEANS > SALINITY/DENSITY > CONDUCTIVITY, EARTH SCIENCE > OCEANS > OCEAN TEMPERATURE > TEMPERATURE PROFILES, EARTH SCIENCE > OCEANS > SALINITY/DENSITY > SALINITY" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:conventions = "CF-1.8, ACDD-1.3" ;
		:id = "PO.DAAC-SMODE-RVCTD" ;
		:uuid = "f8f73c19-7aab-45da-a6b5-d04632077959" ;
		:naming_authority = "gov.nasa" ;
		:featureType = "profile" ;
		:cdm_data_type = "Station" ;
		:source = "TBD" ;
		:platform = "In Situ Ocean-based Platforms > SHIPS > RV Oceanus" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:instrument = "In Situ/Laboratory Instruments > Profilers/Sounders > > > CTD" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:processing_level = "L2" ;
		:standard_name_vocabulary = "CF Standard Name Table v72" ;
		:acknowledgement = "TBD" ;
		:comment = "" ;
		:license = "S-MODE data are considered experimental and not to be used for any purpose for which life or property is potentially at risk. Distributor assumes no responsibility for the manner in which the data are used. Otherwise data are free for public use." ;
		:product_version = "1" ;
		:metadata_link = "https://doi.org/10.5067/SMODE-RVCTD" ;
		:creator_name = "Melissa Omand" ;
		:creator_email = "momand@uri.edu" ;
		:creator_type = "person" ;
		:creator_institution = "URI/" ;
		:institution = "URI/" ;
		:project = "Sub-Mesoscale Ocean Dynamics Experiment (S-MODE)" ;
		:program = "NASA Earth Venture Suborbital-3 (EVS-3)" ;
		:contributor_name = "Frederick Bingham" ;
		:contributor_role = "Project Data Manager" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center, Jet Propulsion Laboratory, NASA" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:sea_name = "Pacific" ;
		:geospatial_lat_min = 16.6695 ;
		:geospatial_lat_max = 16.6695 ;
		:geospatial_lat_units = "degrees" ;
		:geospatial_lat_resolution = "0.1" ;
		:geospatial_lon_min = -146.547666666667 ;
		:geospatial_lon_max = -146.547666666667 ;
		:geospatial_lon_units = "degrees" ;
		:geospatial_lon_resolution = "0.1" ;
		:geospatial_vertical_min = -0.887 ;
		:geospatial_vertical_max = 1053.523 ;
		:geospatial_vertical_resolution = "1" ;
		:geospatial_vertical_units = "m" ;
		:geospatial_vertical_positive = "down" ;
		:time_coverage_start = "16-Aug-2016 20:29:02" ;
		:time_coverage_end = "16-Aug-2016 20:29:02" ;
		:date_created = "01-Sep-2020 14:10:24" ;
}
