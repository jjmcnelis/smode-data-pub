netcdf S-MODE_PFC_waveglider_\#\# {
dimensions:
	upper_time = 90039 ;
	lower_time = 50348 ;
	meteorological_time = 17699 ;
variables:
	double upper_time(upper_time) ;
		upper_time:long_name = "Upper Time of Waveglider measurement" ;
		upper_time:axis = "T" ;
		upper_time:standard_name = "time" ;
		upper_time:units = "days since 1950-01-01T00:00:00" ;
		upper_time:coverage_content_type = "coordinate" ;
	double lower_time(lower_time) ;
		lower_time:long_name = "Lower Time of Waveglider measurement" ;
		lower_time:axis = "T" ;
		lower_time:standard_name = "time" ;
		lower_time:units = "days since 1950-01-01T00:00:00" ;
		lower_time:coverage_content_type = "coordinate" ;
	double upper_longitude(upper_time) ;
		upper_longitude:long_name = "Upper Longitude of Waveglider measurement" ;
		upper_longitude:valid_max = 180. ;
		upper_longitude:valid_min = -180. ;
		upper_longitude:axis = "X" ;
		upper_longitude:standard_name = "longitude" ;
		upper_longitude:units = "degrees_east" ;
		upper_longitude:coverage_content_type = "coordinate" ;
	double lower_longitude(lower_time) ;
		lower_longitude:long_name = "Lower Longitude of Waveglider measurement" ;
		lower_longitude:valid_max = 180. ;
		lower_longitude:valid_min = -180. ;
		lower_longitude:axis = "X" ;
		lower_longitude:standard_name = "longitude" ;
		lower_longitude:units = "degrees_east" ;
		lower_longitude:coverage_content_type = "coordinate" ;
	double upper_latitude(upper_time) ;
		upper_latitude:long_name = "Upper Latitude of Waveglider measurement" ;
		upper_latitude:valid_max = 90. ;
		upper_latitude:valid_min = -90. ;
		upper_latitude:axis = "Y" ;
		upper_latitude:standard_name = "latitude" ;
		upper_latitude:units = "degrees_north" ;
		upper_latitude:coverage_content_type = "coordinate" ;
	double lower_latitude(lower_time) ;
		lower_latitude:_FillValue = NaN ;
		lower_latitude:long_name = "Lower Latitude of Waveglider measurement" ;
		lower_latitude:valid_max = 90. ;
		lower_latitude:valid_min = -90. ;
		lower_latitude:axis = "Y" ;
		lower_latitude:standard_name = "latitude" ;
		lower_latitude:units = "degrees_north" ;
		lower_latitude:coverage_content_type = "coordinate" ;
	double upper_salinity(upper_time) ;
		upper_salinity:_FillValue = NaN ;
		upper_salinity:long_name = "Upper Salinity of Waveglider" ;
		upper_salinity:valid_max = 42. ;
		upper_salinity:valid_min = 2. ;
		upper_salinity:add_offset = 0. ;
		upper_salinity:coorinates = "upper_time upper_latitude upper_longitude" ;
		upper_salinity:scale_factor = 1. ;
		upper_salinity:standard_name = "sea_water_practical_salinity" ;
		upper_salinity:units = "1" ;
		upper_salinity:coverage_content_type = "physicalMeasurement" ;
	double lower_salinity(lower_time) ;
		lower_salinity:_FillValue = NaN ;
		lower_salinity:long_name = "Lower Salinity of Waveglider" ;
		lower_salinity:valid_max = 42. ;
		lower_salinity:valid_min = 2. ;
		lower_salinity:add_offset = 0. ;
		lower_salinity:coorinates = "lower_time lower_latitude lower_longitude" ;
		lower_salinity:scale_factor = 1. ;
		lower_salinity:standard_name = "sea_water_practical_salinity" ;
		lower_salinity:units = "1" ;
		lower_salinity:coverage_content_type = "physicalMeasurement" ;
	double upper_temperature(upper_time) ;
		upper_temperature:_FillValue = NaN ;
		upper_temperature:long_name = "Upper Temperature of Waveglider" ;
		upper_temperature:valid_max = 32. ;
		upper_temperature:valid_min = -1. ;
		upper_temperature:add_offset = 0. ;
		upper_temperature:coorinates = "upper_time upper_latitude upper_longitude" ;
		upper_temperature:scale_factor = 1. ;
		upper_temperature:standard_name = "sea_water_temperature" ;
		upper_temperature:units = "degrees_C" ;
		upper_temperature:coverage_content_type = "physicalMeasurement" ;
	double lower_temperature(lower_time) ;
		lower_temperature:_FillValue = NaN ;
		lower_temperature:long_name = "Lower Temperature of Waveglider" ;
		lower_temperature:valid_max = 32. ;
		lower_temperature:valid_min = -1. ;
		lower_temperature:add_offset = 0. ;
		lower_temperature:coorinates = "lower_time lower_latitude lower_longitude" ;
		lower_temperature:scale_factor = 1. ;
		lower_temperature:standard_name = "sea_water_temperature" ;
		lower_temperature:units = "degrees_C" ;
		lower_temperature:coverage_content_type = "physicalMeasurement" ;
	double upper_pressure(upper_time) ;
		upper_pressure:_FillValue = NaN ;
		upper_pressure:long_name = "Upper Pressure of Waveglider" ;
		upper_pressure:valid_max = 5. ;
		upper_pressure:valid_min = 0. ;
		upper_pressure:add_offset = 0. ;
		upper_pressure:coorinates = "upper_time upper_latitude upper_longitude" ;
		upper_pressure:scale_factor = 1. ;
		upper_pressure:standard_name = "sea_water_pressure" ;
		upper_pressure:units = "dbar" ;
		upper_pressure:coverage_content_type = "physicalMeasurement" ;
	double lower_pressure(lower_time) ;
		lower_pressure:_FillValue = NaN ;
		lower_pressure:long_name = "Lower Pressure of Waveglider" ;
		lower_pressure:valid_max = 10. ;
		lower_pressure:valid_min = 0. ;
		lower_pressure:add_offset = 0. ;
		lower_pressure:coorinates = "lower_time lower_latitude lower_longitude" ;
		lower_pressure:scale_factor = 1. ;
		lower_pressure:standard_name = "sea_water_pressure" ;
		lower_pressure:units = "dbar" ;
		lower_pressure:coverage_content_type = "physicalMeasurement" ;
	double meteorological_time(meteorological_time) ;
		meteorological_time:long_name = "Meteorological Time from an Airmar WX200 instrument on a 1-meter-tall mast" ;
		meteorological_time:axis = "T" ;
		meteorological_time:standard_name = "time" ;
		meteorological_time:units = "days since 1950-01-01T00:00:00" ;
		meteorological_time:coverage_content_type = "coordinate" ;
	double meteorological_longitude(meteorological_time) ;
		meteorological_longitude:_FillValue = NaN ;
		meteorological_longitude:long_name = "Meteorological Longitude from an Airmar WX200 instrument on a 1-meter-tall mast" ;
		meteorological_longitude:valid_max = 180. ;
		meteorological_longitude:valid_min = -180. ;
		meteorological_longitude:axis = "X" ;
		meteorological_longitude:standard_name = "longitude" ;
		meteorological_longitude:units = "degrees_east" ;
		meteorological_longitude:coverage_content_type = "coordinate" ;
	double meteorological_latitude(meteorological_time) ;
		meteorological_latitude:_FillValue = NaN ;
		meteorological_latitude:long_name = "Meteorological Latitude from an Airmar WX200 instrument on a 1-meter-tall mast" ;
		meteorological_latitude:valid_max = 90. ;
		meteorological_latitude:valid_min = -90. ;
		meteorological_latitude:axis = "Y" ;
		meteorological_latitude:standard_name = "latitude" ;
		meteorological_latitude:units = "degrees_north" ;
		meteorological_latitude:coverage_content_type = "coordinate" ;
	double meteorological_wind_direction(meteorological_time) ;
		meteorological_wind_direction:_FillValue = NaN ;
		meteorological_wind_direction:long_name = "Meteorological Wind Direction from an Airmar WX200 instrument on a 1-meter-tall mast" ;
		meteorological_wind_direction:valid_max = 360. ;
		meteorological_wind_direction:valid_min = 0. ;
		meteorological_wind_direction:add_offset = 0. ;
		meteorological_wind_direction:coordinates = "meteorological_time meteorological_latitude meteorological_longitude" ;
		meteorological_wind_direction:scale_factor = 1. ;
		meteorological_wind_direction:standard_name = "wind_from_direction" ;
		meteorological_wind_direction:units = "degree" ;
		meteorological_wind_direction:coverage_content_type = "physicalMeasurement" ;
	double meteorological_wind_speed(meteorological_time) ;
		meteorological_wind_speed:_FillValue = NaN ;
		meteorological_wind_speed:long_name = "Meteorological Wind Speed from an Airmar WX200 instrument on a 1-meter-tall mast" ;
		meteorological_wind_speed:valid_max = 100. ;
		meteorological_wind_speed:valid_min = 0. ;
		meteorological_wind_speed:add_offset = 0. ;
		meteorological_wind_speed:coordinates = "meteorological_time meteorological_latitude meteorological_longitude" ;
		meteorological_wind_speed:scale_factor = 1. ;
		meteorological_wind_speed:standard_name = "wind_speed" ;
		meteorological_wind_speed:units = "knots" ;
		meteorological_wind_speed:coverage_content_type = "physicalMeasurement" ;
	double meteorological_temperature(meteorological_time) ;
		meteorological_temperature:_FillValue = NaN ;
		meteorological_temperature:long_name = "Meteorological Temperature from an Airmar WX200 instrument on a 1-meter-tall mast" ;
		meteorological_temperature:valid_max = 40. ;
		meteorological_temperature:valid_min = 0. ;
		meteorological_temperature:add_offset = 0. ;
		meteorological_temperature:coordinates = "meteorological_time meteorological_latitude meteorological_longitude" ;
		meteorological_temperature:scale_factor = 1. ;
		meteorological_temperature:standard_name = "air_temperature" ;
		meteorological_temperature:units = "degrees_C" ;
		meteorological_temperature:coverage_content_type = "physicalMeasurement" ;
	double meteorological_pressure(meteorological_time) ;
		meteorological_pressure:_FillValue = NaN ;
		meteorological_pressure:long_name = "Meteorological Pressure from an Airmar WX200 instrument on a 1-meter-tall mast" ;
		meteorological_pressure:valid_max = 1030. ;
		meteorological_pressure:valid_min = 900. ;
		meteorological_pressure:add_offset = 0. ;
		meteorological_pressure:coordinates = "meteorological_time meteorological_latitude meteorological_longitude" ;
		meteorological_pressure:scale_factor = 1. ;
		meteorological_pressure:standard_name = "air_pressure" ;
		meteorological_pressure:units = "mbar" ;
		meteorological_pressure:coverage_content_type = "physicalMeasurement" ;

// global attributes:
		:DOI = "10.5067/SMODE-GLID3" ;
		:title = "S-MODE  Pilot Field Campaign Fall 2020 Ocean Temperature and Salinity from Wavegliders<, XXXX>" ;
		:summary = "S-MODE  Pilot Field Campaign Fall 2020 Ocean Temperature and Salinity from Wavegliders<, XXXX>" ;
		:keywords = "EARTH SCIENCE > OCEANS > SALINITY/DENSITY > CONDUCTIVITY, EARTH SCIENCE > OCEANS > OCEAN WINDS > SURFACE WINDS, EARTH SCIENCE > OCEANS > OCEAN TEMPERATURE > TEMPERATURE PROFILES, EARTH SCIENCE > OCEANS > OCEAN CIRCULATION > CURRENT VELOCITY, EARTH SCIENCE > OCEANS > SALINITY/DENSITY > SALINITY, EARTH SCIENCE > OCEANS > OCEAN TEMPERATURE > SURFACE AIR TEMPERATURE, EARTH SCIENCE > OCEANS > OCEAN PRESSURE > SURFACE PRESSURE" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:conventions = "CF-1.8, ACDD-1.3" ;
		:id = "PO.DAAC-SMODE-GLID3" ;
		:uuid = "5a7433df-fc1f-4385-aea9-4b84c6afeea6" ;
		:naming_authority = "gov.nasa" ;
		:featureType = "trajectory" ;
		:cdm_data_type = "Trajectory" ;
		:source = "TBD" ;
		:platform = "In Situ Ocean-based Platforms > USV > WAVEGLIDER" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:instrument = "In Situ/Laboratory Instruments > Recorders/Loggers > > > MMS, In Situ/Laboratory Instruments > Current/Wind Meters > > > CURRENT METERS, In Situ/Laboratory Instruments > Profilers/Sounders > > > CTD" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:processing_level = "L2" ;
		:standard_name_vocabulary = "CF Standard Name Table v72" ;
		:acknowledgement = "TBD" ;
		:comment = "" ;
		:license = "S-MODE data are considered experimental and not to be used for any purpose for which life or property is potentially at risk. Distributor assumes no responsibility for the manner in which the data are used. Otherwise data are free for public use." ;
		:product_version = "1" ;
		:metadata_link = "https://doi.org/10.5067/SMODE-GLID3" ;
		:creator_name = "Tom Farrar" ;
		:creator_email = "jfarrar@whoi.edu" ;
		:creator_type = "person" ;
		:creator_institution = "WHOI/" ;
		:institution = "WHOI/" ;
		:project = "Sub-Mesoscale Ocean Dynamics Experiment (S-MODE)" ;
		:program = "NASA Earth Venture Suborbital-3 (EVS-3)" ;
		:contributor_name = "Frederick Bingham" ;
		:contributor_role = "Project Data Manager" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center, Jet Propulsion Laboratory, NASA" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:sea_name = "Pacific" ;
		:geospatial_lat_min = 9.52764333333333 ;
		:geospatial_lat_max = 13.772675 ;
		:geospatial_lat_units = "degrees" ;
		:geospatial_lat_resolution = "0.1" ;
		:geospatial_lon_min = -126.438033333333 ;
		:geospatial_lon_max = -120.715178333333 ;
		:geospatial_lon_units = "degrees" ;
		:geospatial_lon_resolution = "0.1" ;
		:geospatial_vertical_min = 0.010000229 ;
		:geospatial_vertical_max = 0.40999985 ;
		:geospatial_vertical_resolution = "1" ;
		:geospatial_vertical_units = "m" ;
		:geospatial_vertical_positive = "down" ;
		:time_coverage_start = "24-Aug-2016 00:01:54" ;
		:time_coverage_end = "31-Dec-2016 00:45:51" ;
		:date_created = "01-Sep-2020 14:15:07" ;
}
