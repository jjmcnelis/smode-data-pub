netcdf dopplerscatt-20191206_094944_0422-0474_line09.L2 {
dimensions:
	x = 301 ;
	y = 482 ;
variables:
	double x(x) ;
		x:_FillValue = NaN ;
		x:long_name = "Web Mercator easting" ;
		x:units = "m" ;
		x:valid_min = -1000000. ;
		x:valid_max = 1000000. ;
	double y(y) ;
		y:_FillValue = NaN ;
		y:long_name = "Web Mercator northing" ;
		y:units = "m" ;
		y:valid_min = -1000000. ;
		y:valid_max = 1000000. ;
	double latitude(y) ;
		latitude:_FillValue = NaN ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "Measurement center latitude" ;
		latitude:units = "degrees_north" ;
		latitude:valid_min = -90. ;
		latitude:valid_max = 90. ;
		latitude:coordinates = "spatial_ref" ;
	double longitude(x) ;
		longitude:_FillValue = NaN ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "Measurement center longitude" ;
		longitude:units = "degrees_east" ;
		longitude:valid_min = -180. ;
		longitude:valid_max = 180. ;
		longitude:coordinates = "spatial_ref" ;
	double time(y, x) ;
		time:_FillValue = NaN ;
		time:standard_name = "time" ;
		time:long_name = "Measurement average UTC time." ;
		time:units = "Days after 1950-01-01" ;
		time:valid_min = 0LL ;
		time:valid_max = 36500. ;
		time:grid_mapping = "spatial_ref" ;
		time:coordinates = "spatial_ref" ;
	double wind_speed(y, x) ;
		wind_speed:_FillValue = NaN ;
		wind_speed:description = "m/s" ;
		wind_speed:units = "m s-1" ;
		wind_speed:standard_name = "wind_speed" ;
		wind_speed:long_name = "Neutral wind speed at 10m." ;
		wind_speed:valid_min = 0. ;
		wind_speed:valid_max = 20. ;
		wind_speed:grid_mapping = "spatial_ref" ;
		wind_speed:coordinates = "spatial_ref" ;
	double wind_dir(y, x) ;
		wind_dir:_FillValue = NaN ;
		wind_dir:standard_name = "wind_to_direction" ;
		wind_dir:long_name = "Wind to direction clockwise relative to north." ;
		wind_dir:units = "degrees" ;
		wind_dir:valid_min = -180. ;
		wind_dir:valid_max = 180. ;
		wind_dir:grid_mapping = "spatial_ref" ;
		wind_dir:coordinates = "spatial_ref" ;
	double u_current(y, x) ;
		u_current:_FillValue = NaN ;
		u_current:standard_name = "surface_eastward_sea_water_velocity" ;
		u_current:long_name = "Surface current east component" ;
		u_current:units = "m s-1" ;
		u_current:valid_min = -5. ;
		u_current:valid_max = 5. ;
		u_current:grid_mapping = "spatial_ref" ;
		u_current:coordinates = "spatial_ref" ;
	double v_current(y, x) ;
		v_current:_FillValue = NaN ;
		v_current:standard_name = "surface_northward_sea_water_velocity" ;
		v_current:long_name = "Surface current north component" ;
		v_current:units = "m s-1" ;
		v_current:valid_min = -5. ;
		v_current:valid_max = 5. ;
		v_current:grid_mapping = "spatial_ref" ;
		v_current:coordinates = "spatial_ref" ;
	double u_current_std(y, x) ;
		u_current_std:_FillValue = NaN ;
		u_current_std:long_name = "Surface current east component standard deviation" ;
		u_current_std:units = "m s-1" ;
		u_current_std:valid_min = 0LL ;
		u_current_std:valid_max = 5LL ;
		u_current_std:grid_mapping = "spatial_ref" ;
		u_current_std:coordinates = "spatial_ref" ;
	double v_current_std(y, x) ;
		v_current_std:_FillValue = NaN ;
		v_current_std:long_name = "Surface current north component standard deviation" ;
		v_current_std:units = "m s-1" ;
		v_current_std:valid_min = 0LL ;
		v_current_std:valid_max = 5LL ;
		v_current_std:grid_mapping = "spatial_ref" ;
		v_current_std:coordinates = "spatial_ref" ;
	double tau_x(y, x) ;
		tau_x:_FillValue = NaN ;
		tau_x:description = "m/s" ;
		tau_x:units = "Pa" ;
		tau_x:drag_coefficient = "large-pond-vera" ;
		tau_x:standard_name = "downward_x_stress_at_sea_water_surface" ;
		tau_x:long_name = "Wind stress east component" ;
		tau_x:valid_min = -1. ;
		tau_x:valid_max = 1. ;
		tau_x:grid_mapping = "spatial_ref" ;
		tau_x:coordinates = "spatial_ref" ;
	double tau_y(y, x) ;
		tau_y:_FillValue = NaN ;
		tau_y:description = "m/s" ;
		tau_y:units = "Pa" ;
		tau_y:drag_coefficient = "large-pond-vera" ;
		tau_y:standard_name = "downward_y_stress_at_sea_water_surface" ;
		tau_y:long_name = "Wind stress north component" ;
		tau_y:valid_min = -1. ;
		tau_y:valid_max = 1. ;
		tau_y:grid_mapping = "spatial_ref" ;
		tau_y:coordinates = "spatial_ref" ;
	ubyte flag(y, x) ;
		flag:long_name = "Quality . 1: bad derivatives and smooth data, 2: bad current and winds" ;
		flag:units = "NA" ;
		flag:valid_min = 0LL ;
		flag:valid_max = 255LL ;
		flag:grid_mapping = "spatial_ref" ;
		flag:coordinates = "spatial_ref" ;
	double du_current_dx(y, x) ;
		du_current_dx:_FillValue = NaN ;
		du_current_dx:units = "s-1" ;
		du_current_dx:long_name = "East component of surface current derivative in the east direction" ;
		du_current_dx:valid_min = -0.005 ;
		du_current_dx:valid_max = 0.005 ;
		du_current_dx:grid_mapping = "spatial_ref" ;
		du_current_dx:coordinates = "spatial_ref" ;
	double du_current_dy(y, x) ;
		du_current_dy:_FillValue = NaN ;
		du_current_dy:units = "s-1" ;
		du_current_dy:long_name = "East component of surface current derivative in the north direction" ;
		du_current_dy:valid_min = -0.005 ;
		du_current_dy:valid_max = 0.005 ;
		du_current_dy:grid_mapping = "spatial_ref" ;
		du_current_dy:coordinates = "spatial_ref" ;
	double dv_current_dx(y, x) ;
		dv_current_dx:_FillValue = NaN ;
		dv_current_dx:units = "s-1" ;
		dv_current_dx:long_name = "North component of surface current derivative in the east direction" ;
		dv_current_dx:valid_min = -0.005 ;
		dv_current_dx:valid_max = 0.005 ;
		dv_current_dx:grid_mapping = "spatial_ref" ;
		dv_current_dx:coordinates = "spatial_ref" ;
	double dv_current_dy(y, x) ;
		dv_current_dy:_FillValue = NaN ;
		dv_current_dy:units = "s-1" ;
		dv_current_dy:long_name = "North component of surface current derivative in the north direction" ;
		dv_current_dy:valid_min = -0.005 ;
		dv_current_dy:valid_max = 0.005 ;
		dv_current_dy:grid_mapping = "spatial_ref" ;
		dv_current_dy:coordinates = "spatial_ref" ;
	double surface_current_relative_vorticity(y, x) ;
		surface_current_relative_vorticity:_FillValue = NaN ;
		surface_current_relative_vorticity:units = "s-1" ;
		surface_current_relative_vorticity:long_name = "Surface current relative vorticity" ;
		surface_current_relative_vorticity:valid_min = -0.005 ;
		surface_current_relative_vorticity:valid_max = 0.005 ;
		surface_current_relative_vorticity:grid_mapping = "spatial_ref" ;
		surface_current_relative_vorticity:coordinates = "spatial_ref" ;
	double surface_current_divergence(y, x) ;
		surface_current_divergence:_FillValue = NaN ;
		surface_current_divergence:units = "s-1" ;
		surface_current_divergence:long_name = "Surface current divergence" ;
		surface_current_divergence:valid_min = -0.005 ;
		surface_current_divergence:valid_max = 0.005 ;
		surface_current_divergence:grid_mapping = "spatial_ref" ;
		surface_current_divergence:coordinates = "spatial_ref" ;
	double surface_current_strain_rate(y, x) ;
		surface_current_strain_rate:_FillValue = NaN ;
		surface_current_strain_rate:units = "s-1" ;
		surface_current_strain_rate:long_name = "Surface current strain rate" ;
		surface_current_strain_rate:valid_min = 0LL ;
		surface_current_strain_rate:valid_max = 0.005 ;
		surface_current_strain_rate:grid_mapping = "spatial_ref" ;
		surface_current_strain_rate:coordinates = "spatial_ref" ;
	double du_current_dx_std(y, x) ;
		du_current_dx_std:_FillValue = NaN ;
		du_current_dx_std:units = "s-1" ;
		du_current_dx_std:long_name = "East component of surface current derivative in the east direction standard deviation" ;
		du_current_dx_std:valid_min = 0LL ;
		du_current_dx_std:valid_max = 0.005 ;
		du_current_dx_std:grid_mapping = "spatial_ref" ;
		du_current_dx_std:coordinates = "spatial_ref" ;
	double du_current_dy_std(y, x) ;
		du_current_dy_std:_FillValue = NaN ;
		du_current_dy_std:units = "s-1" ;
		du_current_dy_std:long_name = "East component of surface current derivative in the north direction standard deviation" ;
		du_current_dy_std:valid_min = 0LL ;
		du_current_dy_std:valid_max = 0.005 ;
		du_current_dy_std:grid_mapping = "spatial_ref" ;
		du_current_dy_std:coordinates = "spatial_ref" ;
	double dv_current_dx_std(y, x) ;
		dv_current_dx_std:_FillValue = NaN ;
		dv_current_dx_std:units = "s-1" ;
		dv_current_dx_std:long_name = "North component of surface current derivative in the east direction standard deviation" ;
		dv_current_dx_std:valid_min = 0LL ;
		dv_current_dx_std:valid_max = 0.005 ;
		dv_current_dx_std:grid_mapping = "spatial_ref" ;
		dv_current_dx_std:coordinates = "spatial_ref" ;
	double dv_current_dy_std(y, x) ;
		dv_current_dy_std:_FillValue = NaN ;
		dv_current_dy_std:units = "s-1" ;
		dv_current_dy_std:long_name = "North component of surface current derivative in the north direction standard deviation" ;
		dv_current_dy_std:valid_min = 0LL ;
		dv_current_dy_std:valid_max = 0.005 ;
		dv_current_dy_std:grid_mapping = "spatial_ref" ;
		dv_current_dy_std:coordinates = "spatial_ref" ;
	double surface_current_relative_vorticity_std(y, x) ;
		surface_current_relative_vorticity_std:_FillValue = NaN ;
		surface_current_relative_vorticity_std:units = "s-1" ;
		surface_current_relative_vorticity_std:long_name = "Surface current relative vorticity standard deviation" ;
		surface_current_relative_vorticity_std:valid_min = 0LL ;
		surface_current_relative_vorticity_std:valid_max = 0.005 ;
		surface_current_relative_vorticity_std:grid_mapping = "spatial_ref" ;
		surface_current_relative_vorticity_std:coordinates = "spatial_ref" ;
	double surface_current_divergence_std(y, x) ;
		surface_current_divergence_std:_FillValue = NaN ;
		surface_current_divergence_std:units = "s-1" ;
		surface_current_divergence_std:long_name = "Surface current divergence standard deviation" ;
		surface_current_divergence_std:valid_min = 0LL ;
		surface_current_divergence_std:valid_max = 0.005 ;
		surface_current_divergence_std:grid_mapping = "spatial_ref" ;
		surface_current_divergence_std:coordinates = "spatial_ref" ;
	double dtau_x_dx(y, x) ;
		dtau_x_dx:_FillValue = NaN ;
		dtau_x_dx:units = "N m-3" ;
		dtau_x_dx:long_name = "East component of wind stress derivative in the east direction" ;
		dtau_x_dx:valid_min = -0.0005 ;
		dtau_x_dx:valid_max = 0.0005 ;
		dtau_x_dx:grid_mapping = "spatial_ref" ;
		dtau_x_dx:coordinates = "spatial_ref" ;
	double dtau_x_dy(y, x) ;
		dtau_x_dy:_FillValue = NaN ;
		dtau_x_dy:units = "N m-3" ;
		dtau_x_dy:long_name = "East component of wind stress derivative in the north direction" ;
		dtau_x_dy:valid_min = -0.0005 ;
		dtau_x_dy:valid_max = 0.0005 ;
		dtau_x_dy:grid_mapping = "spatial_ref" ;
		dtau_x_dy:coordinates = "spatial_ref" ;
	double dtau_y_dx(y, x) ;
		dtau_y_dx:_FillValue = NaN ;
		dtau_y_dx:units = "N m-3" ;
		dtau_y_dx:long_name = "North component of wind stress derivative in the east direction" ;
		dtau_y_dx:valid_min = -0.0005 ;
		dtau_y_dx:valid_max = 0.0005 ;
		dtau_y_dx:grid_mapping = "spatial_ref" ;
		dtau_y_dx:coordinates = "spatial_ref" ;
	double dtau_y_dy(y, x) ;
		dtau_y_dy:_FillValue = NaN ;
		dtau_y_dy:units = "N m-3" ;
		dtau_y_dy:long_name = "North component of wind stress derivative in the north direction" ;
		dtau_y_dy:valid_min = -0.0005 ;
		dtau_y_dy:valid_max = 0.0005 ;
		dtau_y_dy:grid_mapping = "spatial_ref" ;
		dtau_y_dy:coordinates = "spatial_ref" ;
	double wind_stress_curl(y, x) ;
		wind_stress_curl:_FillValue = NaN ;
		wind_stress_curl:units = "N m-3" ;
		wind_stress_curl:long_name = "Wind stress curl at the surface" ;
		wind_stress_curl:valid_min = -0.0005 ;
		wind_stress_curl:valid_max = 0.0005 ;
		wind_stress_curl:grid_mapping = "spatial_ref" ;
		wind_stress_curl:coordinates = "spatial_ref" ;
	int64 spatial_ref ;
		spatial_ref:spatial_ref = "PROJCS[\"WGS 84 / Pseudo-Mercator\",GEOGCS[\"WGS 84\",DATUM[\"WGS_1984\",SPHEROID[\"WGS 84\",6378137,298.257223563,AUTHORITY[\"EPSG\",\"7030\"]],AUTHORITY[\"EPSG\",\"6326\"]],PRIMEM[\"Greenwich\",0,AUTHORITY[\"EPSG\",\"8901\"]],UNIT[\"degree\",0.0174532925199433,AUTHORITY[\"EPSG\",\"9122\"]],AUTHORITY[\"EPSG\",\"4326\"]],PROJECTION[\"Mercator_1SP\"],PARAMETER[\"central_meridian\",0],PARAMETER[\"scale_factor\",1],PARAMETER[\"false_easting\",0],PARAMETER[\"false_northing\",0],UNIT[\"metre\",1,AUTHORITY[\"EPSG\",\"9001\"]],AXIS[\"Easting\",EAST],AXIS[\"Northing\",NORTH],EXTENSION[\"PROJ4\",\"+proj=merc +a=6378137 +b=6378137 +lat_ts=0 +lon_0=0 +x_0=0 +y_0=0 +k=1 +units=m +nadgrids=@null +wktext +no_defs\"],AUTHORITY[\"EPSG\",\"3857\"]]" ;
		spatial_ref:crs_wkt = "PROJCS[\"WGS 84 / Pseudo-Mercator\",GEOGCS[\"WGS 84\",DATUM[\"WGS_1984\",SPHEROID[\"WGS 84\",6378137,298.257223563,AUTHORITY[\"EPSG\",\"7030\"]],AUTHORITY[\"EPSG\",\"6326\"]],PRIMEM[\"Greenwich\",0,AUTHORITY[\"EPSG\",\"8901\"]],UNIT[\"degree\",0.0174532925199433,AUTHORITY[\"EPSG\",\"9122\"]],AUTHORITY[\"EPSG\",\"4326\"]],PROJECTION[\"Mercator_1SP\"],PARAMETER[\"central_meridian\",0],PARAMETER[\"scale_factor\",1],PARAMETER[\"false_easting\",0],PARAMETER[\"false_northing\",0],UNIT[\"metre\",1,AUTHORITY[\"EPSG\",\"9001\"]],AXIS[\"Easting\",EAST],AXIS[\"Northing\",NORTH],EXTENSION[\"PROJ4\",\"+proj=merc +a=6378137 +b=6378137 +lat_ts=0 +lon_0=0 +x_0=0 +y_0=0 +k=1 +units=m +nadgrids=@null +wktext +no_defs\"],AUTHORITY[\"EPSG\",\"3857\"]]" ;

// global attributes:
		:cell_size = 400LL ;
		:xmin = -13671142.2768769 ;
		:xmax = -13550895.818709 ;
		:ymin = 4280507.37489517 ;
		:ymax = 4473225.08288703 ;
		:thetamin = 53. ;
		:thetamax = 59. ;
		:xfactormax = "None" ;
		:xfactormin = "None" ;
		:l2a_file_0 = "20191206_094944_0422-0474_line09.L2A.bcolz" ;
		:l2a_file_0_peg_hdg = -28.3527733484922 ;
		:l2a_file_0_peg_lat = 36.5571142180241 ;
		:l2a_file_0_peg_lon = -122.2697756031 ;
		:l2a_file_0_peg_localRadius = 6364290.6188787 ;
		:l2a_file_0_lon0 = -122.2697756031 ;
		:l2a_file_0_lat0 = 36.5571142180241 ;
		:l2a_file_0_grid_spacing = 200. ;
		:l2a_file_0_x_extent = 1000000. ;
		:l2a_file_0_y_extent = 1000000. ;
		:l2a_file_0_projection = "webmercator" ;
		:gl2a_file = "20191206_094944_0422-0474_line09.BDOP.nc" ;
		:line = 9LL ;
		:drag_coefficient = "large-pond-vera" ;
		:title = "DopplerScatt observations from the AITT Field Campaign December 2019" ;
		:summary = "DopplerScatt observations of ocean surface winds currents and from the AITT Field Campaign December 2019" ;
		:creator_name = "E. Rodriguez, A. Wineteer, T. Gal, D. Perkovic-Martin, H. Torres" ;
		:creator_institution = "Jet Propulsion Laboratory, California Institute of Technology" ;
		:creator_email = "ernesto.rodriguez@jpl.nasa.gov" ;
		string :references = "Rodríguez E, Wineteer A, Perkovic-Martin D, Gál T, Stiles BW, Niamsuwan N, Rodriguez Monje R.\nEstimating ocean vector winds and currents using a Ka-band pencil-beam doppler scatterometer.\nRemote Sensing. 2018 Apr;10(4):576." ;
		:feature_type = "grid" ;
		:product_version = "1.0.0" ;
		:date_created = "2020-02-13T22:53:43.261887" ;
		:geospatial_lat_min = "35.85368565113913" ;
		:geospatial_lat_max = "37.24437937456678" ;
		:geospatial_lon_min = "-122.8099605869108" ;
		:geospatial_lon_max = "-121.72976827457576" ;
		:grid_mapping = "spatial_ref" ;
}
