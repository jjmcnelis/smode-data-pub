netcdf S-MODE_PFC_OC2004B_underwayctd_\#\# {
dimensions:
	depth = 69 ;
	time = 259 ;
variables:
	double depth(depth) ;
		depth:_FillValue = NaN ;
		depth:long_name = "Depth of uCTD" ;
		depth:valid_max = 1000. ;
		depth:valid_min = 0. ;
		depth:axis = "Z" ;
		depth:positive = "down" ;
		depth:standard_name = "depth" ;
		depth:units = "m" ;
		depth:coverage_content_type = "coordinate" ;
	double time(time) ;
		time:long_name = "Time of uCTD" ;
		time:axis = "T" ;
		time:standard_name = "time" ;
		time:units = "days since 1950-01-01T00:00:00" ;
		time:coverage_content_type = "coordinate" ;
	double serial_number(time) ;
		serial_number:_FillValue = NaN ;
		serial_number:long_name = "Serial Number of uCTD Probe" ;
		serial_number:coverage_content_type = "referenceInformation" ;
	double latitude(time) ;
		latitude:_FillValue = NaN ;
		latitude:long_name = "Latitude of uCTD" ;
		latitude:valid_max = 90. ;
		latitude:valid_min = -90. ;
		latitude:axis = "Y" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "coordinate" ;
	double longitude(time) ;
		longitude:_FillValue = NaN ;
		longitude:long_name = "Longitude of uCTD" ;
		longitude:valid_max = 180. ;
		longitude:valid_min = -180. ;
		longitude:axis = "X" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "coordinate" ;
	double potential_temperature(time, depth) ;
		potential_temperature:_FillValue = NaN ;
		potential_temperature:long_name = "Potential Temperature of uCTD measurement" ;
		potential_temperature:valid_max = 32. ;
		potential_temperature:valid_min = -1. ;
		potential_temperature:add_offset = 0. ;
		potential_temperature:coordinates = "time depth longitude latitude" ;
		potential_temperature:scale_factor = 1. ;
		potential_temperature:standard_name = "sea_water_potential_temperature" ;
		potential_temperature:units = "degrees_C" ;
		potential_temperature:coverage_content_type = "physicalMeasurement" ;
	double temperature(time, depth) ;
		temperature:_FillValue = NaN ;
		temperature:long_name = "Temperature of uCTD measurement" ;
		temperature:valid_max = 32. ;
		temperature:valid_min = -1. ;
		temperature:add_offset = 0. ;
		temperature:coordinates = "time depth longitude latitude" ;
		temperature:scale_factor = 1. ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "degrees_C" ;
		temperature:coverage_content_type = "physicalMeasurement" ;
	double pressure(time, depth) ;
		pressure:_FillValue = NaN ;
		pressure:long_name = "Pressure of uCTD measurement" ;
		pressure:valid_max = 600. ;
		pressure:valid_min = 0. ;
		pressure:add_offset = 0. ;
		pressure:coordinates = "time depth longitude latitude" ;
		pressure:scale_factor = 1. ;
		pressure:standard_name = "sea_water_pressure" ;
		pressure:units = "dbar" ;
		pressure:coverage_content_type = "physicalMeasurement" ;
	double salinity(time, depth) ;
		salinity:_FillValue = NaN ;
		salinity:long_name = "Salinity of uCTD measurement" ;
		salinity:valid_max = 42. ;
		salinity:valid_min = 2. ;
		salinity:add_offset = 0. ;
		salinity:coordinates = "time depth longitude latitude" ;
		salinity:scale_factor = 1. ;
		salinity:standard_name = "sea_water_practical_salinity" ;
		salinity:units = "1" ;
		salinity:coverage_content_type = "physicalMeasurement" ;
	double eastward_sea_water_velocity(time, depth) ;
		eastward_sea_water_velocity:_FillValue = NaN ;
		eastward_sea_water_velocity:long_name = "Eastward Velocity from ADCP" ;
		eastward_sea_water_velocity:valid_max = 3.11325443716126 ;
		eastward_sea_water_velocity:valid_min = -3.07061233951636 ;
		eastward_sea_water_velocity:add_offset = 0. ;
		eastward_sea_water_velocity:scale_factor = 1. ;
		eastward_sea_water_velocity:standard_name = "eastward_sea_water_velocity" ;
		eastward_sea_water_velocity:units = "m s-1" ;
		eastward_sea_water_velocity:coordinates = "time depth longitude latitude" ;
		eastward_sea_water_velocity:coverage_content_type = "physicalMeasurement" ;
		eastward_sea_water_velocity:comment = "Velocities come from ADCP" ;
	double northward_sea_water_velocity(time, depth) ;
		northward_sea_water_velocity:_FillValue = NaN ;
		northward_sea_water_velocity:long_name = "Northward Velocity from ADCP" ;
		northward_sea_water_velocity:valid_max = 1.98356703246262 ;
		northward_sea_water_velocity:valid_min = -3.05495244808019 ;
		northward_sea_water_velocity:add_offset = 0. ;
		northward_sea_water_velocity:scale_factor = 1. ;
		northward_sea_water_velocity:standard_name = "northward_sea_water_velocity" ;
		northward_sea_water_velocity:units = "m s-1" ;
		northward_sea_water_velocity:coordinates = "time depth longitude latitude" ;
		northward_sea_water_velocity:coverage_content_type = "physicalMeasurement" ;
		northward_sea_water_velocity:comment = "Velocities come from ADCP" ;
	double speed_of_sound_in_sea_water(time, depth) ;
		speed_of_sound_in_sea_water:_FillValue = NaN ;
		speed_of_sound_in_sea_water:long_name = "Speed of Sound in Sea Water of uCTD measurement" ;
		speed_of_sound_in_sea_water:valid_max = 1600. ;
		speed_of_sound_in_sea_water:valid_min = 1400. ;
		speed_of_sound_in_sea_water:add_offset = 0. ;
		speed_of_sound_in_sea_water:coordinates = "time depth longitude latitude" ;
		speed_of_sound_in_sea_water:scale_factor = 1. ;
		speed_of_sound_in_sea_water:standard_name = "speed_of_sound_in_sea_water" ;
		speed_of_sound_in_sea_water:units = "m s-1" ;
		speed_of_sound_in_sea_water:coverage_content_type = "physicalMeasurement" ;
	double sea_water_density(time, depth) ;
		sea_water_density:_FillValue = NaN ;
		sea_water_density:long_name = "Sea Water Density of uCTD measurement" ;
		sea_water_density:valid_max = 30. ;
		sea_water_density:valid_min = 20. ;
		sea_water_density:add_offset = 0. ;
		sea_water_density:coordinates = "time depth longitude latitude" ;
		sea_water_density:scale_factor = 1. ;
		sea_water_density:standard_name = "sea_water_sigma_theta" ;
		sea_water_density:units = "kg m-3" ;
		sea_water_density:coverage_content_type = "physicalMeasurement" ;

// global attributes:
		:DOI = "10.5067/SMODE-RVUCT" ;
		:title = "S-MODE Pilot Field Campaign Fall 2020 Shipboard Underway CTD Measurements R/V Oceanus<, XXXX>" ;
		:summary = "S-MODE Pilot Field Campaign Fall 2020 Shipboard Underway CTD Measurements R/V Oceanus<, XXXX>" ;
		:keywords = "EARTH SCIENCE > OCEANS > SALINITY/DENSITY > CONDUCTIVITY, EARTH SCIENCE > OCEANS > OCEAN TEMPERATURE > TEMPERATURE PROFILES, EARTH SCIENCE > OCEANS > SALINITY/DENSITY > SALINITY" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:conventions = "CF-1.8, ACDD-1.3" ;
		:id = "PO.DAAC-SMODE-RVUCT" ;
		:uuid = "e5cdfd34-eb5f-421a-9576-9fdad6104d13" ;
		:naming_authority = "gov.nasa" ;
		:featureType = "profile" ;
		:cdm_data_type = "Station" ;
		:source = "TBD" ;
		:platform = "In Situ Ocean-based Platforms > SHIPS > RV Oceanus" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:instrument = "In Situ/Laboratory Instruments > Profilers/Sounders > > > CTD" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:processing_level = "L2" ;
		:standard_name_vocabulary = "CF Standard Name Table v72" ;
		:acknowledgement = "TBD" ;
		:comment = "" ;
		:license = "S-MODE data are considered experimental and not to be used for any purpose for which life or property is potentially at risk. Distributor assumes no responsibility for the manner in which the data are used. Otherwise data are free for public use." ;
		:product_version = "1" ;
		:metadata_link = "https://doi.org/10.5067/SMODE-RVUCT" ;
		:creator_name = "Melissa Omand" ;
		:creator_email = "momand@uri.edu" ;
		:creator_type = "person" ;
		:creator_institution = "URI/" ;
		:institution = "URI/" ;
		:project = "Sub-Mesoscale Ocean Dynamics Experiment (S-MODE)" ;
		:program = "NASA Earth Venture Suborbital-3 (EVS-3)" ;
		:contributor_name = "Frederick Bingham" ;
		:contributor_role = "Project Data Manager" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center, Jet Propulsion Laboratory, NASA" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:sea_name = "Pacific" ;
		:geospatial_lat_min = 5.11256141786427 ;
		:geospatial_lat_max = 11.5000350216987 ;
		:geospatial_lat_units = "degrees" ;
		:geospatial_lat_resolution = "0.1" ;
		:geospatial_lon_min = 233.491413283426 ;
		:geospatial_lon_max = 236.499998679269 ;
		:geospatial_lon_units = "degrees" ;
		:geospatial_lon_resolution = "0.1" ;
		:geospatial_vertical_min = 6. ;
		:geospatial_vertical_max = 550. ;
		:geospatial_vertical_resolution = "1" ;
		:geospatial_vertical_units = "m" ;
		:geospatial_vertical_positive = "down" ;
		:time_coverage_start = "21-Aug-2016 21:50:36" ;
		:time_coverage_end = "12-Sep-2016 16:10:21" ;
		:date_created = "01-Sep-2020 14:15:17" ;
}
