9c9
< 		time:units = "days since 1950-01-01T00:00:00" ;
---
> 		time:units = "days since 1950-01-01 00:00:00" ;
12c12
< 		longitude:_FillValue = NaN ;
---
> 		longitude:_FillValue = -9999. ;
16d15
< 		longitude:axis = "X" ;
19c18
< 		longitude:coverage_content_type = "coordinate" ;
---
> 		longitude:coverage_content_type = "referenceInformation" ;
21c20
< 		latitude:_FillValue = NaN ;
---
> 		latitude:_FillValue = -9999. ;
25d23
< 		latitude:axis = "Y" ;
28c26
< 		latitude:coverage_content_type = "coordinate" ;
---
> 		latitude:coverage_content_type = "referenceInformation" ;
30c28
< 		speed_over_ground:_FillValue = NaN ;
---
> 		speed_over_ground:_FillValue = -9999. ;
41c39
< 		course_over_ground:_FillValue = NaN ;
---
> 		course_over_ground:_FillValue = -9999. ;
52c50
< 		pressure_2m:_FillValue = NaN ;
---
> 		pressure_2m:_FillValue = -9999. ;
63c61
< 		pressure_3m:_FillValue = NaN ;
---
> 		pressure_3m:_FillValue = -9999. ;
74c72
< 		density_2m:_FillValue = NaN ;
---
> 		density_2m:_FillValue = -9999. ;
85c83
< 		density_3m:_FillValue = NaN ;
---
> 		density_3m:_FillValue = -9999. ;
96c94
< 		salinity_2m:_FillValue = NaN ;
---
> 		salinity_2m:_FillValue = -9999. ;
107c105
< 		salinity_3m:_FillValue = NaN ;
---
> 		salinity_3m:_FillValue = -9999. ;
118c116
< 		uncorrected_salinity_5m:_FillValue = NaN ;
---
> 		uncorrected_salinity_5m:_FillValue = -9999. ;
129c127
< 		temperature_2m:_FillValue = NaN ;
---
> 		temperature_2m:_FillValue = -9999. ;
140c138
< 		temperature_3m:_FillValue = NaN ;
---
> 		temperature_3m:_FillValue = -9999. ;
151c149
< 		uncorrected_temperature_5m:_FillValue = NaN ;
---
> 		uncorrected_temperature_5m:_FillValue = -9999. ;
162c160
< 		downwelling_longwave_infrared_radiation:_FillValue = NaN ;
---
> 		downwelling_longwave_infrared_radiation:_FillValue = -9999. ;
173c171
< 		downwelling_shortwave_solar_radiation:_FillValue = NaN ;
---
> 		downwelling_shortwave_solar_radiation:_FillValue = -9999. ;
184c182
< 		relative_humidity:_FillValue = NaN ;
---
> 		relative_humidity:_FillValue = -9999. ;
195c193
< 		cumulative_rain:_FillValue = NaN ;
---
> 		cumulative_rain:_FillValue = -9999. ;
206c204
< 		wind_direction:_FillValue = NaN ;
---
> 		wind_direction:_FillValue = -9999. ;
217c215
< 		wind_speed:_FillValue = NaN ;
---
> 		wind_speed:_FillValue = -9999. ;
228c226
< 		ship_heave:_FillValue = NaN ;
---
> 		ship_heave:_FillValue = -9999. ;
239c237
< 		ship_pitch:_FillValue = NaN ;
---
> 		ship_pitch:_FillValue = -9999. ;
250c248
< 		ship_roll:_FillValue = NaN ;
---
> 		ship_roll:_FillValue = -9999. ;
261c259
< 		air_pressure:_FillValue = NaN ;
---
> 		air_pressure:_FillValue = -9999. ;
272c270
< 		air_temperature:_FillValue = NaN ;
---
> 		air_temperature:_FillValue = -9999. ;
290c288
< 		:id = "PO.DAAC-SMODE-RVTSG" ;
---
> 		:id = "PODAAC-SMODE-RVTSG" ;
295c293
< 		:source = "TBD" ;
---
> 		:source = "S-MODE_PFC_OC2004B_thermosalinograph_##.nc.cdl" ;
324,325c322,323
< 		:geospatial_lat_units = "degrees" ;
< 		:geospatial_lat_resolution = "0.1" ;
---
> 		:geospatial_lat_units = "degrees_north" ;
> 		:geospatial_lat_resolution = "0.1 degrees" ;
328,329c326,327
< 		:geospatial_lon_units = "degrees" ;
< 		:geospatial_lon_resolution = "0.1" ;
---
> 		:geospatial_lon_units = "degrees_east" ;
> 		:geospatial_lon_resolution = "0.1 degrees" ;
332,333c330,331
< 		:geospatial_vertical_resolution = "1" ;
< 		:geospatial_vertical_units = "m" ;
---
> 		:geospatial_vertical_resolution = "1 meters" ;
> 		:geospatial_vertical_units = "meters" ;
335,337c333,335
< 		:time_coverage_start = "x" ;
< 		:time_coverage_end = "22-Sep-2016 23:59:55" ;
< 		:date_created = "01-Sep-2020 14:19:07" ;
---
> 		:time_coverage_start = "YYYY-MM-DDTHH:MM:SS" ;
> 		:time_coverage_end = "2016-09-22T23:59:55" ;
> 		:date_created = "2020-09-01T14:19:07" ;
