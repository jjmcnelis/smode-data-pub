10c10
< 		time:units = "days since 1950-01-01T00:00:00" ;
---
> 		time:units = "days since 1950-01-01 00:00:00" ;
13d12
< 		latitude:_FillValue = NaN ;
16,18d14
< 		latitude:valid_max = 90. ;
< 		latitude:valid_min = -90. ;
< 		latitude:axis = "Y" ;
21c17
< 		latitude:coverage_content_type = "coordinate" ;
---
> 		latitude:coverage_content_type = "referenceInformation" ;
23d18
< 		longitude:_FillValue = NaN ;
26,28d20
< 		longitude:valid_max = 180. ;
< 		longitude:valid_min = -180. ;
< 		longitude:axis = "X" ;
31c23
< 		longitude:coverage_content_type = "coordinate" ;
---
> 		longitude:coverage_content_type = "referenceInformation" ;
33c25
< 		speed_over_ground:_FillValue = NaN ;
---
> 		speed_over_ground:_FillValue = -9999. ;
37,38d28
< 		speed_over_ground:add_offset = 0. ;
< 		speed_over_ground:scale_factor = 1. ;
44c34
< 		course_over_ground:_FillValue = NaN ;
---
> 		course_over_ground:_FillValue = -9999. ;
48,49d37
< 		course_over_ground:add_offset = 0. ;
< 		course_over_ground:scale_factor = 1. ;
55c43
< 		heading:_FillValue = NaN ;
---
> 		heading:_FillValue = -9999. ;
59,60d46
< 		heading:add_offset = 0. ;
< 		heading:scale_factor = 1. ;
66c52
< 		eastward_current:_FillValue = NaN ;
---
> 		eastward_current:_FillValue = -9999. ;
70,71d55
< 		eastward_current:add_offset = 0. ;
< 		eastward_current:scale_factor = 1. ;
77c61
< 		northward_current:_FillValue = NaN ;
---
> 		northward_current:_FillValue = -9999. ;
81,82d64
< 		northward_current:add_offset = 0. ;
< 		northward_current:scale_factor = 1. ;
88c70
< 		wind_speed_relative_to_earth_18m:_FillValue = NaN ;
---
> 		wind_speed_relative_to_earth_18m:_FillValue = -9999. ;
92,93d73
< 		wind_speed_relative_to_earth_18m:add_offset = 0. ;
< 		wind_speed_relative_to_earth_18m:scale_factor = 1. ;
99c79
< 		wind_direction_relative_to_earth:_FillValue = NaN ;
---
> 		wind_direction_relative_to_earth:_FillValue = -9999. ;
103,104d82
< 		wind_direction_relative_to_earth:add_offset = 0. ;
< 		wind_direction_relative_to_earth:scale_factor = 1. ;
110c88
< 		wind_speed_relative_to_earth:_FillValue = NaN ;
---
> 		wind_speed_relative_to_earth:_FillValue = -9999. ;
114,115d91
< 		wind_speed_relative_to_earth:add_offset = 0. ;
< 		wind_speed_relative_to_earth:scale_factor = 1. ;
121c97
< 		neutral_wind_speed_relative_to_earth:_FillValue = NaN ;
---
> 		neutral_wind_speed_relative_to_earth:_FillValue = -9999. ;
125,126d100
< 		neutral_wind_speed_relative_to_earth:add_offset = 0. ;
< 		neutral_wind_speed_relative_to_earth:scale_factor = 1. ;
132c106
< 		wind_speed_relative_to_water_18m:_FillValue = NaN ;
---
> 		wind_speed_relative_to_water_18m:_FillValue = -9999. ;
136,137d109
< 		wind_speed_relative_to_water_18m:add_offset = 0. ;
< 		wind_speed_relative_to_water_18m:scale_factor = 1. ;
143c115
< 		wind_direction_relative_to_water:_FillValue = NaN ;
---
> 		wind_direction_relative_to_water:_FillValue = -9999. ;
147,148d118
< 		wind_direction_relative_to_water:add_offset = 0. ;
< 		wind_direction_relative_to_water:scale_factor = 1. ;
154c124
< 		wind_speed_relative_to_water_2m:_FillValue = NaN ;
---
> 		wind_speed_relative_to_water_2m:_FillValue = -9999. ;
158,159d127
< 		wind_speed_relative_to_water_2m:add_offset = 0. ;
< 		wind_speed_relative_to_water_2m:scale_factor = 1. ;
165c133
< 		wind_speed_relative_to_water_10m:_FillValue = NaN ;
---
> 		wind_speed_relative_to_water_10m:_FillValue = -9999. ;
169,170d136
< 		wind_speed_relative_to_water_10m:add_offset = 0. ;
< 		wind_speed_relative_to_water_10m:scale_factor = 1. ;
176c142
< 		neutral_wind_speed_relative_to_water:_FillValue = NaN ;
---
> 		neutral_wind_speed_relative_to_water:_FillValue = -9999. ;
180,181d145
< 		neutral_wind_speed_relative_to_water:add_offset = 0. ;
< 		neutral_wind_speed_relative_to_water:scale_factor = 1. ;
187c151
< 		air_temperature_16p5m:_FillValue = NaN ;
---
> 		air_temperature_16p5m:_FillValue = -9999. ;
192,193d155
< 		air_temperature_16p5m:add_offset = 0. ;
< 		air_temperature_16p5m:scale_factor = 1. ;
199c161
< 		air_temperature:_FillValue = NaN ;
---
> 		air_temperature:_FillValue = -9999. ;
204,205d165
< 		air_temperature:add_offset = 0. ;
< 		air_temperature:scale_factor = 1. ;
211c171
< 		near_sea_surface_temperature_5cm:_FillValue = NaN ;
---
> 		near_sea_surface_temperature_5cm:_FillValue = -9999. ;
215,216d174
< 		near_sea_surface_temperature_5cm:add_offset = 0. ;
< 		near_sea_surface_temperature_5cm:scale_factor = 1. ;
222c180
< 		near_sea_surface_temperature_2m:_FillValue = NaN ;
---
> 		near_sea_surface_temperature_2m:_FillValue = -9999. ;
226,227d183
< 		near_sea_surface_temperature_2m:add_offset = 0. ;
< 		near_sea_surface_temperature_2m:scale_factor = 1. ;
233c189
< 		near_sea_surface_temperature_3m:_FillValue = NaN ;
---
> 		near_sea_surface_temperature_3m:_FillValue = -9999. ;
237,238d192
< 		near_sea_surface_temperature_3m:add_offset = 0. ;
< 		near_sea_surface_temperature_3m:scale_factor = 1. ;
244c198
< 		near_sea_surface_temperature_5m:_FillValue = NaN ;
---
> 		near_sea_surface_temperature_5m:_FillValue = -9999. ;
248,249d201
< 		near_sea_surface_temperature_5m:add_offset = 0. ;
< 		near_sea_surface_temperature_5m:scale_factor = 1. ;
255c207
< 		relative_humidity_16p5m:_FillValue = NaN ;
---
> 		relative_humidity_16p5m:_FillValue = -9999. ;
260,261d211
< 		relative_humidity_16p5m:add_offset = 0. ;
< 		relative_humidity_16p5m:scale_factor = 1. ;
263c213
< 		relative_humidity_16p5m:units = "%" ;
---
> 		relative_humidity_16p5m:units = "1" ;
267c217
< 		relative_humidity_2m:_FillValue = NaN ;
---
> 		relative_humidity_2m:_FillValue = -9999. ;
272,273d221
< 		relative_humidity_2m:add_offset = 0. ;
< 		relative_humidity_2m:scale_factor = 1. ;
275c223
< 		relative_humidity_2m:units = "%" ;
---
> 		relative_humidity_2m:units = "1" ;
279c227
< 		relative_humidity_10m:_FillValue = NaN ;
---
> 		relative_humidity_10m:_FillValue = -9999. ;
284,285d231
< 		relative_humidity_10m:add_offset = 0. ;
< 		relative_humidity_10m:scale_factor = 1. ;
287c233
< 		relative_humidity_10m:units = "%" ;
---
> 		relative_humidity_10m:units = "1" ;
291c237
< 		pressure:_FillValue = NaN ;
---
> 		pressure:_FillValue = -9999. ;
295,296d240
< 		pressure:add_offset = 0. ;
< 		pressure:scale_factor = 1. ;
302c246
< 		specific_humidity_16p5m:_FillValue = NaN ;
---
> 		specific_humidity_16p5m:_FillValue = -9999. ;
307,308d250
< 		specific_humidity_16p5m:add_offset = 0. ;
< 		specific_humidity_16p5m:scale_factor = 1. ;
314c256
< 		specific_humidity_2m:_FillValue = NaN ;
---
> 		specific_humidity_2m:_FillValue = -9999. ;
319,320d260
< 		specific_humidity_2m:add_offset = 0. ;
< 		specific_humidity_2m:scale_factor = 1. ;
326c266
< 		specific_humidity_10m:_FillValue = NaN ;
---
> 		specific_humidity_10m:_FillValue = -9999. ;
331,332d270
< 		specific_humidity_10m:add_offset = 0. ;
< 		specific_humidity_10m:scale_factor = 1. ;
338c276
< 		specific_humidity_sea_surface:_FillValue = NaN ;
---
> 		specific_humidity_sea_surface:_FillValue = -9999. ;
343,344d280
< 		specific_humidity_sea_surface:add_offset = 0. ;
< 		specific_humidity_sea_surface:scale_factor = 1. ;
350c286
< 		sss:_FillValue = NaN ;
---
> 		sss:_FillValue = -9999. ;
354,355d289
< 		sss:add_offset = 0. ;
< 		sss:scale_factor = 1. ;
357a292
> 		sss:comments = "SSS is assumed to be a ratio because of units=1. Provide more details about physical units in this field, e.g. (cm3 cm-3)" ;
361c296
< 		salinity_2m:_FillValue = NaN ;
---
> 		salinity_2m:_FillValue = -9999. ;
365,366d299
< 		salinity_2m:add_offset = 0. ;
< 		salinity_2m:scale_factor = 1. ;
372c305
< 		salinity_3m:_FillValue = NaN ;
---
> 		salinity_3m:_FillValue = -9999. ;
376,377d308
< 		salinity_3m:add_offset = 0. ;
< 		salinity_3m:scale_factor = 1. ;
383c314
< 		salinity_5m:_FillValue = NaN ;
---
> 		salinity_5m:_FillValue = -9999. ;
387,388d317
< 		salinity_5m:add_offset = 0. ;
< 		salinity_5m:scale_factor = 1. ;
394c323
< 		precipitation_rate:_FillValue = NaN ;
---
> 		precipitation_rate:_FillValue = -9999. ;
398,399d326
< 		precipitation_rate:add_offset = 0. ;
< 		precipitation_rate:scale_factor = 1. ;
405c332
< 		evaporation_rate:_FillValue = NaN ;
---
> 		evaporation_rate:_FillValue = -9999. ;
409,410d335
< 		evaporation_rate:add_offset = 0. ;
< 		evaporation_rate:scale_factor = 1. ;
423c348
< 		:id = "PO.DAAC-SMODE-RVMET" ;
---
> 		:id = "PODAAC-SMODE-RVMET" ;
428c353
< 		:source = "TBD" ;
---
> 		:source = "S-MODE_PFC_OC2004B_meteorology_##.nc.cdl" ;
457,458c382,383
< 		:geospatial_lat_units = "degrees" ;
< 		:geospatial_lat_resolution = "0.1" ;
---
> 		:geospatial_lat_units = "degrees_north" ;
> 		:geospatial_lat_resolution = "0.1 degrees" ;
461,462c386,387
< 		:geospatial_lon_units = "degrees" ;
< 		:geospatial_lon_resolution = "0.1" ;
---
> 		:geospatial_lon_units = "degrees_east" ;
> 		:geospatial_lon_resolution = "0.1 degrees" ;
465,466c390,391
< 		:geospatial_vertical_resolution = "1" ;
< 		:geospatial_vertical_units = "m" ;
---
> 		:geospatial_vertical_resolution = "1 meters" ;
> 		:geospatial_vertical_units = "meters" ;
468,470c393,395
< 		:time_coverage_start = "20-Aug-2016 00:00:30" ;
< 		:time_coverage_end = "18-Sep-2016 23:59:30" ;
< 		:date_created = "01-Sep-2020 14:11:36" ;
---
> 		:time_coverage_start = "2016-08-20T00:00:30" ;
> 		:time_coverage_end = "2016-09-18T23:59:30" ;
> 		:date_created = "2020-09-01T14:11:36" ;
