netcdf S-MODE_PFC_OC2004B_adcp_\#\# {
dimensions:
	time = 18593 ;
	depth = 60 ;
	trajectory = 1 ;
variables:
	double trajectory(trajectory) ;
		trajectory:standard_name = "trajectory" ;
		trajectory:cf_role = "trajectory_id" ;
	double time(time) ;
		time:long_name = "Time of ADCP measurement" ;
		time:axis = "T" ;
		time:standard_name = "time" ;
		time:units = "days since 1950-01-01 00:00:00" ;
		time:coverage_content_type = "coordinate" ;
	double depth(time, depth) ;
		depth:long_name = "Depth of ADCP measurement" ;
		depth:valid_max = 1000. ;
		depth:valid_min = 0. ;
		depth:axis = "Z" ;
		depth:positive = "down" ;
		depth:standard_name = "depth" ;
		depth:units = "m" ;
		depth:coverage_content_type = "coordinate" ;
	double longitude(time) ;
		longitude:long_name = "Longitude of ADCP measurement" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "referenceInformation" ;
	double latitude(time) ;
		latitude:long_name = "Latitude of ADCP measurement" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "referenceInformation" ;
	double zonal_velocity_component(time, depth) ;
		zonal_velocity_component:_FillValue = -9999. ;
		zonal_velocity_component:long_name = "Zonal velocity component of ADCP measurement" ;
		zonal_velocity_component:valid_max = 5. ;
		zonal_velocity_component:valid_min = -5. ;
		zonal_velocity_component:coordinates = "time latitude longitude depth trajectory" ;
		zonal_velocity_component:standard_name = "seawater_x_velocity" ;
		zonal_velocity_component:units = "m s-1" ;
		zonal_velocity_component:coverage_content_type = "physicalMeasurement" ;
	double meridional_velocity_component(time, depth) ;
		meridional_velocity_component:_FillValue = -9999. ;
		meridional_velocity_component:long_name = "Meridional velocity component of ADCP measurement" ;
		meridional_velocity_component:valid_max = 5. ;
		meridional_velocity_component:valid_min = -5. ;
		meridional_velocity_component:coordinates = "time latitude longitude depth trajectory" ;
		meridional_velocity_component:standard_name = "seawater_y_velocity" ;
		meridional_velocity_component:units = "m s-1" ;
		meridional_velocity_component:coverage_content_type = "physicalMeasurement" ;
	double ship_speed(time) ;
		ship_speed:_FillValue = -9999. ;
		ship_speed:long_name = "Ship zonal velocity component during ADCP measurement" ;
		ship_speed:valid_max = 20. ;
		ship_speed:valid_min = 0. ;
		ship_speed:coordinates = "time latitude longitude depth" ;
		ship_speed:standard_name = "platform_speed_wrt_ground" ;
		ship_speed:units = "m s-1" ;
		ship_speed:coverage_content_type = "physicalMeasurement" ;
	double ship_direction(time) ;
		ship_direction:_FillValue = -9999. ;
		ship_direction:long_name = "Direction of ship during ADCP measurement" ;
		ship_direction:valid_max = 180. ;
		ship_direction:valid_min = -180. ;
		ship_direction:coordinates = "time latitude longitude depth trajectory" ;
		ship_direction:standard_name = "ship_dir" ;
		ship_direction:units = "degrees" ;
		ship_direction:comment = "Ship directions are expressed in degrees normal" ;
		ship_direction:coverage_content_type = "physicalMeasurement" ;
	double amplitude(time, depth) ;
		amplitude:_FillValue = -9999. ;
		amplitude:long_name = "Received signal strength of ADCP measurement" ;
		amplitude:valid_max = 212. ;
		amplitude:valid_min = 12. ;
		amplitude:coordinates = "time latitude longitude depth trajectory" ;
		amplitude:standard_name = "signal_strength" ;
		amplitude:coverage_content_type = "physicalMeasurement" ;
	double percent_good(time, depth) ;
		percent_good:_FillValue = -9999. ;
		percent_good:long_name = "Percent of good pings of ADCP measurement" ;
		percent_good:valid_max = 100. ;
		percent_good:valid_min = 0. ;
		percent_good:coordinates = "time latitude longitude depth trajectory" ;
		percent_good:standard_name = "percent of good pings" ;
		percent_good:coverage_content_type = "physicalMeasurement" ;
	double status_flag(time, depth) ;
		status_flag:_FillValue = -9999. ;
		status_flag:long_name = "Editing flags of ADCP measurement" ;
		status_flag:missing_value = -1. ;
		status_flag:valid_max = 7. ;
		status_flag:valid_min = 0. ;
		status_flag:flag_values = 0., 1., 2., 3., 4., 5., 6., 7. ;
		status_flag:flag_meanings = "good bin_bad percent_good_bad bin_and_percent_good_bad range_bad range_and_bin_bad range_and_percent_good_bad range_and_percent_good_and_bin_bad" ;
		status_flag:standard_name = "status_flag" ;
		status_flag:coordinates = "time latitude longitude depth trajectory" ;
		status_flag:coverage_content_type = "referenceInformation" ;
		status_flag:comment = "Zero indicates good data. For more information see: https://currents.soest.hawaii.edu/docs/adcp_doc/pflags_doc/" ;
	double temperature(time) ;
		temperature:_FillValue = -9999. ;
		temperature:long_name = "Temperature of ADCP transducer" ;
		temperature:valid_max = 32. ;
		temperature:valid_min = -1. ;
		temperature:coordinates = "time latitude longitude depth trajectory" ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "degrees_C" ;
		temperature:coverage_content_type = "physicalMeasurement" ;
}
