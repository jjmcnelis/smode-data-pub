netcdf S-MODE_PFC_surfacedrifter_\#\# {
dimensions:
	time = 48 ;
	trajectory = 1 ;
variables:
	int trajectory(trajectory) ;
        trajectory:long_name = "Unique identifier for each feature instance" ;
        trajectory:cf_role = "trajectory_id" ;
	double time(trajectory, time) ;
		time:long_name = "Time of Salinity Drifter measurement" ;
		time:axis = "T" ;
		time:standard_name = "time" ;
		time:units = "days since 1950-01-01 00:00:00" ;
		time:coverage_content_type = "coordinate" ;
	double longitude(trajectory, time) ;
		longitude:_FillValue = -9999. ;
		longitude:long_name = "Longitude of Salinity Drifter measurement" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "referenceInformation" ;
	double latitude(trajectory, time) ;
		longitude:_FillValue = -9999. ;
		latitude:long_name = "Latitude of Salinity Drifter measurement" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "referenceInformation" ;
	double temperature_18cm(trajectory, time) ;
		temperature_18cm:_FillValue = -9999. ;
		temperature_18cm:long_name = "Sea water temperature at 18cm" ;
		temperature_18cm:valid_max = 32. ;
		temperature_18cm:valid_min = -1. ;
		temperature_18cm:coordinates = "time latitude longitude" ;
		temperature_18cm:standard_name = "sea_water_temperature" ;
		temperature_18cm:units = "degrees_C" ;
		temperature_18cm:coverage_content_type = "physicalMeasurement" ;
		temperature_18cm:comment = "Notice that T(18-cm)  is a hull-sensor that is sensitive to inside-hull temperature. In particular, during the first half hour , these temperatures are not correct." ;
	double temperature_36cm(trajectory, time) ;
		temperature_36cm:_FillValue = -9999. ;
		temperature_36cm:long_name = "Sea water temperature at 36cm" ;
		temperature_36cm:valid_max = 32. ;
		temperature_36cm:valid_min = -1. ;
		temperature_36cm:coordinates = "time latitude longitude" ;
		temperature_36cm:standard_name = "sea_water_temperature" ;
		temperature_36cm:units = "degrees_C" ;
		temperature_36cm:coverage_content_type = "physicalMeasurement" ;
	double salinity_36cm(trajectory, time) ;
		salinity_36cm:_FillValue = -9999. ;
		salinity_36cm:long_name = "Sea water salinity at 36cm" ;
		salinity_36cm:valid_max = 42. ;
		salinity_36cm:valid_min = 2. ;
		salinity_36cm:coordinates = "time latitude longitude" ;
		salinity_36cm:standard_name = "sea_water_practical_salinity" ;
		salinity_36cm:units = "1" ;
		salinity_36cm:comments = "Salinity is assumed to be a ratio because of units=1. Provide more details about physical units in this field, e.g. (cm3 cm-3) for volumetric ratio." ;	
		salinity_36cm:coverage_content_type = "physicalMeasurement" ;

// global attributes:
		:DOI = "10.5067/SMODE-DRIFT" ;
		:title = "S-MODE  Pilot Field Campaign Fall 2020 Position Data from Surface Drifters<, XXXX>" ;
		:summary = "S-MODE  Pilot Field Campaign Fall 2020 Position Data from Surface Drifters<, XXXX>" ;
		:keywords = "EARTH SCIENCE > OCEANS > OCEAN TEMPERATURE > TEMPERATURE PROFILES, EARTH SCIENCE > OCEANS > SALINITY/DENSITY > SALINITY" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:conventions = "CF-1.8, ACDD-1.3" ;
		:id = "PODAAC-SMODE-DRIFT" ;
		:uuid = "9094f9a1-80d7-4b59-b79d-2303d9860d6a" ;
		:naming_authority = "gov.nasa" ;
		:featureType = "trajectory" ;
		:cdm_data_type = "Trajectory" ;
		:source = "S-MODE_PFC_surfacedrifter_\#\#.nc" ;
		:platform = "In Situ Ocean-based Platforms > BUOYS > BUOYS" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:instrument = "In Situ/Laboratory Instruments > Current/Wind Meters > > > DRIFTING BUOYS" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:processing_level = "L2" ;
		:standard_name_vocabulary = "CF Standard Name Table v72" ;
		:acknowledgement = "TBD" ;
		:comment = "" ;
		:license = "S-MODE data are considered experimental and not to be used for any purpose for which life or property is potentially at risk. Distributor assumes no responsibility for the manner in which the data are used. Otherwise data are free for public use." ;
		:product_version = "1" ;
		:metadata_link = "https://doi.org/10.5067/SMODE-DRIFT" ;
		:creator_name = "Andrey Shcherbina" ;
		:creator_email = "shcher@uw.edu" ;
		:creator_type = "person" ;
		:creator_institution = "UWA/" ;
		:institution = "UWA/" ;
		:project = "Sub-Mesoscale Ocean Dynamics Experiment (S-MODE)" ;
		:program = "NASA Earth Venture Suborbital-3 (EVS-3)" ;
		:contributor_name = "Frederick Bingham" ;
		:contributor_role = "Project Data Manager" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center, Jet Propulsion Laboratory, NASA" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:sea_name = "Pacific" ;
		:geospatial_lat_min = 10.5048 ;
		:geospatial_lat_max = 10.5094 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = "0.1 degrees" ;
		:geospatial_lon_min = -124.1476 ;
		:geospatial_lon_max = -124.138 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = "0.1 degrees" ;
		:geospatial_vertical_min = 0.18 ;
		:geospatial_vertical_max = 0.36 ;
		:geospatial_vertical_resolution = "1 meters" ;
		:geospatial_vertical_units = "meters" ;
		:geospatial_vertical_positive = "down" ;
		:time_coverage_start = "2017-11-09T13:10:10" ;
		:time_coverage_end = "2017-11-09T17:05:10" ;
		:date_created = "2020-09-01T14:19:24" ;
}
