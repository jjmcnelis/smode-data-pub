netcdf S-MODE_PFC_slocumglider_\#\# {
dimensions:
	time = 1615 ;
	profile = 46 ;
variables:
	int profile(profile) ;
        profile:long_name = "Unique identifier for each feature instance" ;
        profile:cf_role = "profile_id" ;
	double latitude(time) ;
		longitude:_FillValue = NaN ;
		latitude:long_name = "Latitude" ;
		latitude:valid_max = 90. ;
		latitude:valid_min = -90. ;
		latitude:axis = "Y" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "referenceInformation" ;
	double longitude(time) ;
		longitude:_FillValue = NaN ;
		longitude:long_name = "Longitude" ;
		longitude:valid_max = 180. ;
		longitude:valid_min = -180. ;
		longitude:axis = "X" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "referenceInformation" ;
	double time(time) ;
		sample_time:long_name = "Time" ;
		sample_time:axis = "T" ;
		sample_time:standard_name = "time" ;
		sample_time:units = "days since 1950-01-01 00:00:00" ;
		sample_time:coverage_content_type = "coordinate" ;
	double temperature(time) ;
		temperature:_FillValue = NaN ;
		temperature:long_name = "Temperature" ;
		temperature:valid_max = 32. ;
		temperature:valid_min = -1. ;
		temperature:add_offset = 0. ;
		temperature:coordinates = "time latitude longitude" ;
		temperature:scale_factor = 1. ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "degrees_C" ;
		temperature:coverage_content_type = "physicalMeasurement" ;
		temperature:comment = "corrected for first-order lag" ;
	double original_temperature(time) ;
		original_temperature:_FillValue = NaN ;
		original_temperature:long_name = "Original Sci Reported Temperature" ;
		original_temperature:valid_max = 32. ;
		original_temperature:valid_min = -1. ;
		original_temperature:add_offset = 0. ;
		original_temperature:coordinates = "time latitude longitude" ;
		original_temperature:scale_factor = 1. ;
		original_temperature:standard_name = "sea_water_temperature" ;
		original_temperature:units = "degrees_C" ;
		original_temperature:coverage_content_type = "physicalMeasurement" ;
	double conductivity(time) ;
		conductivity:_FillValue = NaN ;
		conductivity:long_name = "Conductivity" ;
		conductivity:valid_max = 60. ;
		conductivity:valid_min = 0. ;
		conductivity:add_offset = 0. ;
		conductivity:coordinates = "time latitude longitude" ;
		conductivity:scale_factor = 1. ;
		conductivity:standard_name = "sea_water_electrical_conductivity" ;
		conductivity:units = "S m-1" ;
		conductivity:coverage_content_type = "physicalMeasurement" ;
		conductivity:comment = "corrected for first-order lag" ;
	double original_conductivity(time) ;
		original_conductivity:_FillValue = NaN ;
		original_conductivity:long_name = "Original Sci Reported Conductivity" ;
		original_conductivity:valid_max = 60. ;
		original_conductivity:valid_min = 0. ;
		original_conductivity:add_offset = 0. ;
		original_conductivity:coordinates = "time latitude longitude" ;
		original_conductivity:scale_factor = 1. ;
		original_conductivity:standard_name = "sea_water_electrical_conductivity" ;
		original_conductivity:units = "S m-1" ;
		original_conductivity:coverage_content_type = "physicalMeasurement" ;
		original_conductivity:comment = "corrected for first-order lag" ;
	double salinity(time) ;
		salinity:_FillValue = NaN ;
		salinity:long_name = "Salinity" ;
		salinity:valid_max = 42. ;
		salinity:valid_min = 2. ;
		salinity:add_offset = 0. ;
		salinity:coordinates = "time latitude longitude" ;
		salinity:scale_factor = 1. ;
		salinity:standard_name = "sea_water_practical_salinity" ;
		salinity:units = "1" ;
		salinity:coverage_content_type = "physicalMeasurement" ;
	double depth(time) ;
		depth:_FillValue = NaN ;
		depth:long_name = "Depth" ;
		depth:valid_max = 1500. ;
		depth:valid_min = 0. ;
		depth:axis = "Z" ;
		depth:positive = "down" ;
		depth:standard_name = "depth" ;
		depth:units = "m" ;
		depth:coverage_content_type = "coordinate" ;
	double profile_start_index(profile_number) ;
		profile_start_index:coverage_content_type = "referenceInformation" ;
	double profile_end_index(profile_number) ;
		profile_end_index:coverage_content_type = "referenceInformation" ;
	double temperature_flag(time) ;
		temperature_flag:_FillValue = NaN ;
		temperature_flag:long_name = "Temperature editing flags" ;
		temperature_flag:missing_value = -1. ;
		temperature_flag:valid_max = 9. ;
		temperature_flag:valid_min = 1. ;
		temperature_flag:flag_values = 1., 2., 4., 5., 6., 9. ;
		temperature_flag:flag_meanings = "1: Good; 2: Range tests, Bad; 4: Digit Rollover, Spike tests, Density Inversion Probably Bad; 5:  Shallow/Deep Gradient, Pressure Gap, Probably Bad; 6: Increasing Pressure, Bad; 9: No QC Performed" ;
		temperature_flag:add_offset = 0. ;
		temperature_flag:scale_factor = 1. ;
		temperature_flag:standard_name = "status_flag" ;
		temperature_flag:coordinates = "depth time latitude longitude" ;
		temperature_flag:coverage_content_type = "referenceInformation" ;
		temperature_flag:comment = "One indicates good data." ;
	double salt_flag(time) ;
		salt_flag:_FillValue = NaN ;
		salt_flag:long_name = "Salinity editing flags" ;
		salt_flag:missing_value = -1. ;
		salt_flag:valid_max = 9. ;
		salt_flag:valid_min = 1. ;
		salt_flag:flag_values = 0., 1., 2., 3., 4., 5., 6., 7. ;
		salt_flag:flag_meanings = "1: Good; 2: Range tests, Bad; 4: Digit Rollover, Spike tests, Density Inversion Probably Bad; 5:  Shallow/Deep Gradient, Pressure Gap, Probably Bad; 6: Increasing Pressure, Bad; 9: No QC Performed" ;
		salt_flag:add_offset = 0. ;
		salt_flag:scale_factor = 1. ;
		salt_flag:standard_name = "status_flag" ;
		salt_flag:coordinates = "depth time latitude longitude" ;
		salt_flag:coverage_content_type = "referenceInformation" ;
		salt_flag:comment = "Zero indicates good data." ;

// global attributes:
		:DOI = "10.5067/SMODE-GLID2" ;
		:title = "S-MODE  Pilot Field Campaign Fall 2020 Temperature and Salinity from Slocum Gliders<, XXXX>" ;
		:summary = "S-MODE  Pilot Field Campaign Fall 2020 Temperature and Salinity from Slocum Gliders<, XXXX>" ;
		:keywords = "EARTH SCIENCE > OCEANS > SALINITY/DENSITY > CONDUCTIVITY, EARTH SCIENCE > OCEANS > OCEAN TEMPERATURE > TEMPERATURE PROFILES, EARTH SCIENCE > OCEANS > SALINITY/DENSITY > SALINITY" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:conventions = "CF-1.8, ACDD-1.3" ;
		:id = "PO.DAAC-SMODE-GLID2" ;
		:uuid = "4c6ea1a7-1c96-4746-8a81-e58480b5ff3a" ;
		:naming_authority = "gov.nasa" ;
		:featureType = "trajectoryProfile" ;
		:cdm_data_type = "TrajectoryProfile" ;
		:source = "TBD" ;
		:platform = "In Situ Ocean-based Platforms > USV" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:instrument = "In Situ/Laboratory Instruments > Profilers/Sounders > > > CTD" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:processing_level = "L3" ;
		:standard_name_vocabulary = "CF Standard Name Table v73" ;
		:acknowledgement = "TBD" ;
		:comment = "" ;
		:license = "S-MODE data are considered experimental and not to be used for any purpose for which life or property is potentially at risk. Distributor assumes no responsibility for the manner in which the data are used. Otherwise data are free for public use." ;
		:product_version = "2" ;
		:metadata_link = "https://doi.org/10.5067/SMODE-GLID2" ;
		:creator_name = "Joseph D\'Addezio" ;
		:creator_email = "joseph.daddezio@nrlssc.navy.mil" ;
		:creator_type = "person" ;
		:creator_institution = "NRL/" ;
		:institution = "NRL/" ;
		:project = "Sub-Mesoscale Ocean Dynamics Experiment (S-MODE)" ;
		:program = "NASA Earth Venture Suborbital-3 (EVS-3)" ;
		:contributor_name = "Frederick Bingham" ;
		:contributor_role = "Project Data Manager" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center, Jet Propulsion Laboratory, NASA" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:sea_name = "Pacific" ;
		:geospatial_lat_min = 39.23934f ;
		:geospatial_lat_max = 39.26562f ;
		:geospatial_lat_units = "degrees" ;
		:geospatial_lat_resolution = "0.1" ;
		:geospatial_lon_min = -74.21561f ;
		:geospatial_lon_max = -74.20511f ;
		:geospatial_lon_units = "degrees" ;
		:geospatial_lon_resolution = "0.1" ;
		:geospatial_vertical_min = 0.2077447f ;
		:geospatial_vertical_max = 64.09405f ;
		:geospatial_vertical_resolution = "1" ;
		:geospatial_vertical_units = "m" ;
		:geospatial_vertical_positive = "down" ;
		:time_coverage_start = "27-Aug-6662" ;
		:time_coverage_end = "27-Dec-6697" ;
		:date_created = "01-Sep-2020 16:37:30" ;
}
