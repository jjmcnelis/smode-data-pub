netcdf S-MODE_PFC_saildrone_\#\# {
dimensions:
	time = 4609 ;
variables:
	double time(time) ;
		time:long_name = "Time of Saildrone" ;
		time:axis = "T" ;
		time:standard_name = "time" ;
		time:units = "days since 1950-01-01T00:00:00" ;
		time:coverage_content_type = "coordinate" ;
	double longitude(time) ;
		longitude:_FillValue = NaN ;
		longitude:long_name = "Longitude of Saildrone" ;
		longitude:valid_max = 180. ;
		longitude:valid_min = -180. ;
		longitude:axis = "X" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "coordinate" ;
	double latitude(time) ;
		latitude:_FillValue = NaN ;
		latitude:long_name = "Latitude of Saildrone" ;
		latitude:valid_max = 90. ;
		latitude:valid_min = -90. ;
		latitude:axis = "Y" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "coordinate" ;
	double sst(time) ;
		sst:_FillValue = NaN ;
		sst:long_name = "Sea Surface Temperature" ;
		sst:valid_max = 32. ;
		sst:valid_min = -1. ;
		sst:add_offset = 0. ;
		sst:scale_factor = 1. ;
		sst:standard_name = "sea_surface_temperature" ;
		sst:units = "degrees_C" ;
		sst:coordinates = "time latitude longitude" ;
		sst:coverage_content_type = "physicalMeasurement" ;
	double sss(time) ;
		sss:_FillValue = NaN ;
		sss:long_name = "Sea Surface Salinity" ;
		sss:valid_max = 42. ;
		sss:valid_min = 2. ;
		sss:add_offset = 0. ;
		sss:scale_factor = 1. ;
		sss:standard_name = "sea_water_practical_salinity" ;
		sss:units = "1" ;
		sss:coordinates = "time latitude longitude" ;
		sss:coverage_content_type = "physicalMeasurement" ;
	double solar_radiation(time) ;
		solar_radiation:_FillValue = NaN ;
		solar_radiation:long_name = "Solar Radiation" ;
		solar_radiation:valid_max = 1500. ;
		solar_radiation:valid_min = 0. ;
		solar_radiation:add_offset = 0. ;
		solar_radiation:scale_factor = 1. ;
		solar_radiation:standard_name = "downwelling_shortwave_flux_in_air" ;
		solar_radiation:units = "W m-2" ;
		solar_radiation:coordinates = "time latitude longitude" ;
		solar_radiation:coverage_content_type = "physicalMeasurement" ;
	double long_radiation(time) ;
		long_radiation:_FillValue = NaN ;
		long_radiation:long_name = "Longwave Radiation" ;
		long_radiation:valid_max = 600. ;
		long_radiation:valid_min = 0. ;
		long_radiation:add_offset = 0. ;
		long_radiation:scale_factor = 1. ;
		long_radiation:standard_name = "surface_upwelling_longwave_flux_in_air" ;
		long_radiation:units = "W m-2" ;
		long_radiation:coordinates = "time latitude longitude" ;
		long_radiation:coverage_content_type = "physicalMeasurement" ;
	double pressure(time) ;
		pressure:_FillValue = NaN ;
		pressure:long_name = "Sea Level Pressure" ;
		pressure:valid_max = 1020. ;
		pressure:valid_min = 1000. ;
		pressure:add_offset = 0. ;
		pressure:scale_factor = 1. ;
		pressure:standard_name = "air_pressure_at_sea_level" ;
		pressure:units = "hPa" ;
		pressure:coordinates = "time latitude longitude" ;
		pressure:coverage_content_type = "physicalMeasurement" ;
	double wind_direction(time) ;
		wind_direction:_FillValue = NaN ;
		wind_direction:long_name = "Wind Direction" ;
		wind_direction:valid_max = 180. ;
		wind_direction:valid_min = -180. ;
		wind_direction:add_offset = 0. ;
		wind_direction:scale_factor = 1. ;
		wind_direction:standard_name = "wind_to_direction" ;
		wind_direction:units = "degrees" ;
		wind_direction:coordinates = "time latitude longitude" ;
		wind_direction:coverage_content_type = "physicalMeasurement" ;
		wind_direction:comment = "Angle increases clockwise. 0deg is southerly; 90deg westerly; -90deg easterly; 180deg northerly" ;
	double wind_speed_5m(time) ;
		wind_speed_5m:_FillValue = NaN ;
		wind_speed_5m:long_name = "Wind Speed at 5m" ;
		wind_speed_5m:valid_max = 11.986 ;
		wind_speed_5m:valid_min = 0. ;
		wind_speed_5m:add_offset = 0. ;
		wind_speed_5m:scale_factor = 1. ;
		wind_speed_5m:standard_name = "wind_speed" ;
		wind_speed_5m:units = "m s-1" ;
		wind_speed_5m:coordinates = "time latitude longitude" ;
		wind_speed_5m:coverage_content_type = "physicalMeasurement" ;
	double relative_humidity_2m(time) ;
		relative_humidity_2m:_FillValue = NaN ;
		relative_humidity_2m:long_name = "Relative Humidity at 2.4m" ;
		relative_humidity_2m:valid_max = 100. ;
		relative_humidity_2m:valid_min = 0. ;
		relative_humidity_2m:add_offset = 0. ;
		relative_humidity_2m:scale_factor = 1. ;
		relative_humidity_2m:standard_name = "relative_humidity" ;
		relative_humidity_2m:units = "%" ;
		relative_humidity_2m:coordinates = "time latitude longitude" ;
		relative_humidity_2m:coverage_content_type = "physicalMeasurement" ;
	double specific_humidity_2m(time) ;
		specific_humidity_2m:_FillValue = NaN ;
		specific_humidity_2m:long_name = "Specific Humidity at 2.4m" ;
		specific_humidity_2m:valid_max = 21.185 ;
		specific_humidity_2m:valid_min = 16.274 ;
		specific_humidity_2m:add_offset = 0. ;
		specific_humidity_2m:scale_factor = 1. ;
		specific_humidity_2m:standard_name = "specific_humidity" ;
		specific_humidity_2m:units = "g kg-1" ;
		specific_humidity_2m:coordinates = "time latitude longitude" ;
		specific_humidity_2m:coverage_content_type = "physicalMeasurement" ;
	double air_temperature_2m(time) ;
		air_temperature_2m:_FillValue = NaN ;
		air_temperature_2m:long_name = "Air Temperature at 2.4m" ;
		air_temperature_2m:valid_max = 28.343 ;
		air_temperature_2m:valid_min = 23.316 ;
		air_temperature_2m:add_offset = 0. ;
		air_temperature_2m:scale_factor = 1. ;
		air_temperature_2m:standard_name = "air_temperature" ;
		air_temperature_2m:units = "degrees_C" ;
		air_temperature_2m:coordinates = "time latitude longitude" ;
		air_temperature_2m:coverage_content_type = "physicalMeasurement" ;
	double wind_speed_10m(time) ;
		wind_speed_10m:_FillValue = NaN ;
		wind_speed_10m:long_name = "Wind Speed at 10m" ;
		wind_speed_10m:valid_max = 12.811 ;
		wind_speed_10m:valid_min = 0. ;
		wind_speed_10m:add_offset = 0. ;
		wind_speed_10m:scale_factor = 1. ;
		wind_speed_10m:standard_name = "wind_speed" ;
		wind_speed_10m:units = "m s-1" ;
		wind_speed_10m:coordinates = "time latitude longitude" ;
		wind_speed_10m:coverage_content_type = "physicalMeasurement" ;
	double relative_humidity_10m(time) ;
		relative_humidity_10m:_FillValue = NaN ;
		relative_humidity_10m:long_name = "Relative Humidity at 10m" ;
		relative_humidity_10m:valid_max = 100. ;
		relative_humidity_10m:valid_min = 0. ;
		relative_humidity_10m:add_offset = 0. ;
		relative_humidity_10m:scale_factor = 1. ;
		relative_humidity_10m:standard_name = "relative_humidity" ;
		relative_humidity_10m:units = "%" ;
		relative_humidity_10m:coordinates = "time latitude longitude" ;
		relative_humidity_10m:coverage_content_type = "physicalMeasurement" ;
	double specific_humidity_10m(time) ;
		specific_humidity_10m:_FillValue = NaN ;
		specific_humidity_10m:long_name = "Specific Humidity at 10m" ;
		specific_humidity_10m:valid_max = 20.932 ;
		specific_humidity_10m:valid_min = 15.958 ;
		specific_humidity_10m:add_offset = 0. ;
		specific_humidity_10m:scale_factor = 1. ;
		specific_humidity_10m:standard_name = "specific_humidity" ;
		specific_humidity_10m:units = "g kg-1" ;
		specific_humidity_10m:coordinates = "time latitude longitude" ;
		specific_humidity_10m:coverage_content_type = "physicalMeasurement" ;
	double air_temperature_10m(time) ;
		air_temperature_10m:_FillValue = NaN ;
		air_temperature_10m:long_name = "Air Temperature at 10m" ;
		air_temperature_10m:valid_max = 28.302 ;
		air_temperature_10m:valid_min = 22.878 ;
		air_temperature_10m:add_offset = 0. ;
		air_temperature_10m:scale_factor = 1. ;
		air_temperature_10m:standard_name = "air_temperature" ;
		air_temperature_10m:units = "degrees_C" ;
		air_temperature_10m:coordinates = "time latitude longitude" ;
		air_temperature_10m:coverage_content_type = "physicalMeasurement" ;

// global attributes:
		:DOI = "10.5067/SMODE-SDRON" ;
		:title = "S-MODE  Pilot Field Campaign Fall 2020 Temperature and Salinity from Saildrones<, XXXX>" ;
		:summary = "S-MODE  Pilot Field Campaign Fall 2020 Temperature and Salinity from Saildrones<, XXXX>" ;
		:keywords = "EARTH SCIENCE > ATMOSPHERE > OCEAN WINDS > SURFACE WINDS, EARTH SCIENCE > OCEANS > SALINITY/DENSITY > CONDUCTIVITY, EARTH SCIENCE > OCEANS > OCEAN OPTICS > CHLOROPHYLL, EARTH SCIENCE > OCEANS > SALINITY/DENSITY > SALINITY, EARTH SCIENCE > OCEANS > OCEAN TEMPERATURE > SEA SURFACE TEMPERATURE, EARTH SCIENCE > ATMOSPHERE > ATMOSPHERIC PRESSURE > ATMOSPHERIC PRESSURE MEASUREMENTS, EARTH SCIENCE > ATMOSPHERE > ATMOSPHERIC TEMPERATURE > AIR TEMPERATURE, EARTH SCIENCE > OCEANS > OCEAN CHEMISTRY > OXYGEN" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:conventions = "CF-1.8, ACDD-1.3" ;
		:id = "PO.DAAC-SMODE-SDRON" ;
		:uuid = "344d2690-234f-44d4-b1af-8d464bc725bc" ;
		:naming_authority = "gov.nasa" ;
		:featureType = "trajectory" ;
		:cdm_data_type = "Trajectory" ;
		:source = "TBD" ;
		:platform = "In Situ Ocean-based Platforms > USV > Saildrone" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:instrument = "In Situ/Laboratory Instruments > Profilers/Sounders > Acoustic Sounders > > ADCP" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:processing_level = "L2" ;
		:standard_name_vocabulary = "CF Standard Name Table v72" ;
		:acknowledgement = "TBD" ;
		:comment = "" ;
		:license = "S-MODE data are considered experimental and not to be used for any purpose for which life or property is potentially at risk. Distributor assumes no responsibility for the manner in which the data are used. Otherwise data are free for public use." ;
		:product_version = "1" ;
		:metadata_link = "https://doi.org/10.5067/SMODE-SDRON" ;
		:creator_name = "Cesar B Rocha" ;
		:creator_email = "crocha@whoi.edu" ;
		:creator_type = "person" ;
		:creator_institution = "WHOI/" ;
		:institution = "WHOI/" ;
		:project = "Sub-Mesoscale Ocean Dynamics Experiment (S-MODE)" ;
		:program = "NASA Earth Venture Suborbital-3 (EVS-3)" ;
		:contributor_name = "Frederick Bingham" ;
		:contributor_role = "Project Data Manager" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center, Jet Propulsion Laboratory, NASA" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:sea_name = "Pacific" ;
		:geospatial_lat_min = 10.88961448 ;
		:geospatial_lat_max = 10.88961448 ;
		:geospatial_lat_units = "degrees" ;
		:geospatial_lat_resolution = "0.1" ;
		:geospatial_lon_min = -125.08657088 ;
		:geospatial_lon_max = -124.54938688 ;
		:geospatial_lon_units = "degrees" ;
		:geospatial_lon_resolution = "0.1" ;
		:geospatial_vertical_min = 1006.1575 ;
		:geospatial_vertical_max = 1015.41 ;
		:geospatial_vertical_resolution = "1" ;
		:geospatial_vertical_units = "m" ;
		:geospatial_vertical_positive = "down" ;
		:time_coverage_start = "16-Oct-2017" ;
		:time_coverage_end = "17-Nov-2017" ;
		:date_created = "01-Sep-2020 14:13:03" ;
}
