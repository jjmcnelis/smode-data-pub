netcdf S-MODE_PFC_lagrangianfloat_\#\# {
dimensions:
	ctd_time = 343588 ;
	depth = 2 ;
	fast_time = 8897670 ;
	gps_time = 1808 ;
variables:
	double ctd_depth(depth, ctd_time) ;
		ctd_depth:_FillValue = NaN ;
		ctd_depth:instrument = "2 Sea-Bird Scientific SBE 41 CTD units at top and bottom of float" ;
		ctd_depth:long_name = "Depth at the two CTD units" ;
		ctd_depth:valid_max = 200., 200. ;
		ctd_depth:valid_min = 0., 0. ;
		ctd_depth:axis = "Z" ;
		ctd_depth:positive = "down" ;
		ctd_depth:standard_name = "depth" ;
		ctd_depth:units = "m" ;
		ctd_depth:coverage_content_type = "coordinate" ;
	double float_depth(ctd_time) ;
		float_depth:_FillValue = NaN ;
		float_depth:instrument = "2 Sea-Bird Scientific SBE 41 CTD units at top and bottom of float" ;
		float_depth:long_name = "Depth at the float center" ;
		float_depth:valid_max = 200. ;
		float_depth:valid_min = 0. ;
		float_depth:axis = "Z" ;
		float_depth:positive = "down" ;
		float_depth:standard_name = "depth" ;
		float_depth:units = "m" ;
		float_depth:coverage_content_type = "coordinate" ;
	double fast_depth(fast_time) ;
		fast_depth:_FillValue = NaN ;
		fast_depth:instrument = "Druck PDCR 910-200" ;
		fast_depth:long_name = "Depth at the float center" ;
		fast_depth:valid_max = 200. ;
		fast_depth:valid_min = 0. ;
		fast_depth:axis = "Z" ;
		fast_depth:positive = "down" ;
		fast_depth:standard_name = "depth" ;
		fast_depth:units = "m" ;
		fast_depth:coverage_content_type = "coordinate" ;
	double time(gps_time) ;
		time:instrument = "GARMIN GPS 15H/L" ;
		time:long_name = "Time of GARMIN GPS 15H/L" ;
		time:axis = "T" ;
		time:standard_name = "time" ;
		time:units = "days since 1950-01-01T00:00:00" ;
		time:coverage_content_type = "coordinate" ;
	double longitude(gps_time) ;
		longitude:_FillValue = NaN ;
		longitude:instrument = "GARMIN GPS 15H/L" ;
		longitude:long_name = "Longitude of GARMIN GPS 15H/L" ;
		longitude:valid_max = 180. ;
		longitude:valid_min = -180. ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "coordinate" ;
		longitude:axis = "Y" ;
	double latitude(gps_time) ;
		latitude:_FillValue = NaN ;
		latitude:instrument = "GARMIN GPS 15H/L" ;
		latitude:long_name = "Latitude of GARMIN GPS 15H/L" ;
		latitude:valid_max = 90. ;
		latitude:valid_min = -90. ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "coordinate" ;
	double ctd_time(ctd_time) ;
		ctd_time:instrument = "2 Sea-Bird Scientific SBE 41 CTD units at top and bottom of float" ;
		ctd_time:long_name = "Time of Sea-Bird Scientific SBE 41" ;
		ctd_time:axis = "T" ;
		ctd_time:standard_name = "time" ;
		ctd_time:units = "days since 1950-01-01T00:00:00" ;
		ctd_time:coverage_content_type = "coordinate" ;
	double ctd_temperature(depth, ctd_time) ;
		ctd_temperature:_FillValue = NaN ;
		ctd_temperature:instrument = "2 Sea-Bird Scientific SBE 41 CTD units at top and bottom of float" ;
		ctd_temperature:long_name = "Sea Water Temperature at the two CTD units" ;
		ctd_temperature:valid_max = 32. ;
		ctd_temperature:valid_min = -1. ;
		ctd_temperature:add_offset = 0. ;
		ctd_temperature:scale_factor = 1. ;
		ctd_temperature:standard_name = "sea_water_temperature" ;
		ctd_temperature:units = "degrees_C" ;
		ctd_temperature:coordinates = "ctd_time ctd_depth" ;
		ctd_temperature:coverage_content_type = "physicalMeasurement" ;
	double ctd_salinity(depth, ctd_time) ;
		ctd_salinity:_FillValue = NaN ;
		ctd_salinity:instrument = "2 Sea-Bird Scientific SBE 41 CTD units at top and bottom of float" ;
		ctd_salinity:long_name = "Sea Water Practical Salinity at the two CTD units" ;
		ctd_salinity:valid_max = 42. ;
		ctd_salinity:valid_min = 2. ;
		ctd_salinity:add_offset = 0. ;
		ctd_salinity:scale_factor = 1. ;
		ctd_salinity:standard_name = "sea_water_practical_salinity" ;
		ctd_salinity:units = "1" ;
		ctd_salinity:coordinates = "ctd_time ctd_depth" ;
		ctd_salinity:coverage_content_type = "physicalMeasurement" ;
	double float_pressure(ctd_time) ;
		float_pressure:_FillValue = NaN ;
		float_pressure:instrument = "2 Sea-Bird Scientific SBE 41 CTD units at top and bottom of float" ;
		float_pressure:long_name = "Pressure at the float center" ;
		float_pressure:valid_max = 200. ;
		float_pressure:valid_min = 0. ;
		float_pressure:add_offset = 0. ;
		float_pressure:scale_factor = 1. ;
		float_pressure:standard_name = "sea_water_pressure" ;
		float_pressure:units = "dbar" ;
		float_pressure:coordinates = "ctd_time ctd_depth" ;
		float_pressure:coverage_content_type = "physicalMeasurement" ;
	double ctd_pressure(depth, ctd_time) ;
		ctd_pressure:_FillValue = NaN ;
		ctd_pressure:instrument = "2 Sea-Bird Scientific SBE 41 CTD units at top and bottom of float" ;
		ctd_pressure:long_name = "Pressure at the two CTD units" ;
		ctd_pressure:valid_max = 200. ;
		ctd_pressure:valid_min = 0. ;
		ctd_pressure:add_offset = 0. ;
		ctd_pressure:scale_factor = 1. ;
		ctd_pressure:standard_name = "sea_water_pressure" ;
		ctd_pressure:units = "dbar" ;
		ctd_pressure:coordinates = "ctd_time ctd_depth" ;
		ctd_pressure:coverage_content_type = "physicalMeasurement" ;
	double fast_time(fast_time) ;
		fast_time:instrument = "Druck PDCR 910-200" ;
		fast_time:long_name = "Time of Druck PDCR 910-200" ;
		fast_time:axis = "T" ;
		fast_time:standard_name = "time" ;
		fast_time:units = "days since 1950-01-01T00:00:00" ;
		fast_time:coverage_content_type = "coordinate" ;
	double fast_pressure(fast_time) ;
		fast_pressure:_FillValue = NaN ;
		fast_pressure:instrument = "Druck PDCR 910-200" ;
		fast_pressure:long_name = "Fast Pressure at the float center" ;
		fast_pressure:valid_max = 200. ;
		fast_pressure:valid_min = 0. ;
		fast_pressure:add_offset = 0. ;
		fast_pressure:scale_factor = 1. ;
		fast_pressure:standard_name = "sea_water_pressure" ;
		fast_pressure:units = "dbar" ;
		fast_pressure:coordinates = "ctd_time ctd_depth" ;
		fast_pressure:coverage_content_type = "physicalMeasurement" ;

// global attributes:
		:DOI = "10.5067/SMODE-FLOAT" ;
		:title = "S-MODE  Pilot Field Campaign Fall 2020 Ocean Temperature and Salinity from Lagrangian Floats<, XXXX>" ;
		:summary = "S-MODE  Pilot Field Campaign Fall 2020 Ocean Temperature and Salinity from Lagrangian Floats<, XXXX>" ;
		:keywords = "EARTH SCIENCE > OCEANS > SALINITY/DENSITY > CONDUCTIVITY, EARTH SCIENCE > OCEANS > SALINITY/DENSITY > SALINITY, EARTH SCIENCE > OCEANS > OCEAN TEMPERATURE > TEMPERATURE PROFILES" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:conventions = "CF-1.8, ACDD-1.3" ;
		:id = "PO.DAAC-SMODE-FLOAT" ;
		:uuid = "ca63b056-e895-4723-9fb2-fc2fedc66c01" ;
		:naming_authority = "gov.nasa" ;
		:featureType = "timeSeries" ;
		:cdm_data_type = "Trajectory" ;
		:source = "TBD" ;
		:platform = "In Situ Ocean-based Platforms > FLOATS >" ;
		:platform_vocabulary = "GCMD platform keywords" ;
		:instrument = "In Situ/Laboratory Instruments > Profilers/Sounders > > > CTD" ;
		:instrument_vocabulary = "GCMD instrument keywords" ;
		:processing_level = "L2" ;
		:standard_name_vocabulary = "CF Standard Name Table v72" ;
		:acknowledgement = "TBD" ;
		:comment = "" ;
		:license = "S-MODE data are considered experimental and not to be used for any purpose for which life or property is potentially at risk. Distributor assumes no responsibility for the manner in which the data are used. Otherwise data are free for public use." ;
		:product_version = "1" ;
		:metadata_link = "https://doi.org/10.5067/SMODE-FLOAT" ;
		:creator_name = "Andrey Shcherbina" ;
		:creator_email = "shcher@uw.edu" ;
		:creator_type = "person" ;
		:creator_institution = "UWA/" ;
		:institution = "UWA/" ;
		:project = "Sub-Mesoscale Ocean Dynamics Experiment (S-MODE)" ;
		:program = "NASA Earth Venture Suborbital-3 (EVS-3)" ;
		:contributor_name = "Frederick Bingham" ;
		:contributor_role = "Project Data Manager" ;
		:publisher_name = "Physical Oceanography Distributed Active Archive Center, Jet Propulsion Laboratory, NASA" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:sea_name = "Pacific" ;
		:geospatial_lat_min = 7.85503149032593 ;
		:geospatial_lat_max = 11.8912620544434 ;
		:geospatial_lat_units = "degrees" ;
		:geospatial_lat_resolution = "0.1" ;
		:geospatial_lon_min = -125.015312194824 ;
		:geospatial_lon_max = -108.951736450195 ;
		:geospatial_lon_units = "degrees" ;
		:geospatial_lon_resolution = "0.1" ;
		:geospatial_vertical_min = 9.02827726415439e-05 ;
		:geospatial_vertical_max = 160.111795419475 ;
		:geospatial_vertical_resolution = "1" ;
		:geospatial_vertical_units = "m" ;
		:geospatial_vertical_positive = "down" ;
		:time_coverage_start = "26-Aug-2016 18:38:07" ;
		:time_coverage_end = "12-Dec-2016 13:18:19" ;
		:date_created = "01-Sep-2020 14:11:19" ;
}
